//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccLz.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccLz_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccLz_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccLz(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccLz_rom Thresholding_Batch_0_Thresholding_BatccLz_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccvx.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccvx_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccvx_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccvx(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccvx_rom Thresholding_Batch_0_Thresholding_Batccvx_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbAo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcbAo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbAo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcbAo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcbAo_rom Thresholding_Batch_0_Thresholding_BatcbAo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActCeG.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActCeG_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActCeG_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActCeG(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActCeG_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActCeG_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/hdl/finn_design_wrapper.v

//Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
//--------------------------------------------------------------------------------
//Tool Version: Vivado v.2020.1.1 (lin64) Build 2960000 Wed Aug  5 22:57:21 MDT 2020
//Date        : Sat Jan 30 13:23:55 2021
//Host        : finn_dev_grgov running 64-bit unknown
//Command     : generate_target finn_design_wrapper.bd
//Design      : finn_design_wrapper
//Purpose     : IP block netlist
//--------------------------------------------------------------------------------
`timescale 1 ps / 1 ps

module finn_design_wrapper
   (ap_clk,
    ap_rst_n,
    m_axis_0_tdata,
    m_axis_0_tready,
    m_axis_0_tvalid,
    m_axis_1_tdata,
    m_axis_1_tready,
    m_axis_1_tvalid,
    m_axis_2_tdata,
    m_axis_2_tready,
    m_axis_2_tvalid,
    s_axis_0_tdata,
    s_axis_0_tready,
    s_axis_0_tvalid,
    s_axis_1_tdata,
    s_axis_1_tready,
    s_axis_1_tvalid,
    s_axis_2_tdata,
    s_axis_2_tready,
    s_axis_2_tvalid);
  input ap_clk;
  input ap_rst_n;
  output [7:0]m_axis_0_tdata;
  input m_axis_0_tready;
  output m_axis_0_tvalid;
  output [7:0]m_axis_1_tdata;
  input m_axis_1_tready;
  output m_axis_1_tvalid;
  output [7:0]m_axis_2_tdata;
  input m_axis_2_tready;
  output m_axis_2_tvalid;
  input [7:0]s_axis_0_tdata;
  output s_axis_0_tready;
  input s_axis_0_tvalid;
  input [7:0]s_axis_1_tdata;
  output s_axis_1_tready;
  input s_axis_1_tvalid;
  input [15:0]s_axis_2_tdata;
  output s_axis_2_tready;
  input s_axis_2_tvalid;

  wire ap_clk;
  wire ap_rst_n;
  wire [7:0]m_axis_0_tdata;
  wire m_axis_0_tready;
  wire m_axis_0_tvalid;
  wire [7:0]m_axis_1_tdata;
  wire m_axis_1_tready;
  wire m_axis_1_tvalid;
  wire [7:0]m_axis_2_tdata;
  wire m_axis_2_tready;
  wire m_axis_2_tvalid;
  wire [7:0]s_axis_0_tdata;
  wire s_axis_0_tready;
  wire s_axis_0_tvalid;
  wire [7:0]s_axis_1_tdata;
  wire s_axis_1_tready;
  wire s_axis_1_tvalid;
  wire [15:0]s_axis_2_tdata;
  wire s_axis_2_tready;
  wire s_axis_2_tvalid;

  finn_design finn_design_i
       (.ap_clk(ap_clk),
        .ap_rst_n(ap_rst_n),
        .m_axis_0_tdata(m_axis_0_tdata),
        .m_axis_0_tready(m_axis_0_tready),
        .m_axis_0_tvalid(m_axis_0_tvalid),
        .m_axis_1_tdata(m_axis_1_tdata),
        .m_axis_1_tready(m_axis_1_tready),
        .m_axis_1_tvalid(m_axis_1_tvalid),
        .m_axis_2_tdata(m_axis_2_tdata),
        .m_axis_2_tready(m_axis_2_tready),
        .m_axis_2_tvalid(m_axis_2_tvalid),
        .s_axis_0_tdata(s_axis_0_tdata),
        .s_axis_0_tready(s_axis_0_tready),
        .s_axis_0_tvalid(s_axis_0_tvalid),
        .s_axis_1_tdata(s_axis_1_tdata),
        .s_axis_1_tready(s_axis_1_tready),
        .s_axis_1_tvalid(s_axis_1_tvalid),
        .s_axis_2_tdata(s_axis_2_tdata),
        .s_axis_2_tready(s_axis_2_tready),
        .s_axis_2_tvalid(s_axis_2_tvalid));
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/e911/StreamingFIFO_4.v


module StreamingFIFO_4(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [95:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [95:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(96)
)
StreamingFIFO_4_StreamingFIFO_4
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_StreamingFCLayer_6jw.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

(* use_dsp = "no" *) module StreamingFCLayer_Batch_4_StreamingFCLayer_6jw_Mul_LUT_0(a, b, p);
input[4 - 1 : 0] a; 
input[4 - 1 : 0] b; 
output[8 - 1 : 0] p;

assign p = $signed(a) * $signed(b);
endmodule
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_StreamingFCLayer_6jw(
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



StreamingFCLayer_Batch_4_StreamingFCLayer_6jw_Mul_LUT_0 StreamingFCLayer_Batch_4_StreamingFCLayer_6jw_Mul_LUT_0_U(
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbyn.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbyn_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbyn_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbyn(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbyn_rom Thresholding_Batch_0_Thresholding_Batcbyn_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actyd2.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actyd2_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actyd2_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actyd2(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actyd2_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actyd2_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/bc91/hdl/verilog/StreamingFCLayer_Batch_6_Matrix_Vector_Activa.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingFCLayer_Batch_6_Matrix_Vector_Activa (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY,
        weight_V_V_TDATA,
        weight_V_V_TVALID,
        weight_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [7:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;
input  [7:0] weight_V_V_TDATA;
input   weight_V_V_TVALID;
output   weight_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;
reg weight_V_V_TREADY;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln248_fu_2165_p2;
wire   [0:0] icmp_ln252_fu_2180_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln289_reg_6766;
reg    weight_V_V_TDATA_blk_n;
reg   [10:0] i_0_reg_1625;
reg    ap_predicate_op540_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [10:0] i_fu_2171_p2;
wire   [7:0] inElem_V_1_fu_2961_p258;
wire   [7:0] trunc_ln321_fu_3479_p1;
wire   [0:0] icmp_ln271_fu_4766_p2;
reg   [0:0] icmp_ln271_reg_6751;
wire   [3:0] trunc_ln647_fu_4772_p1;
reg  signed [3:0] trunc_ln647_reg_6756;
reg  signed [3:0] p_Result_s_reg_6761;
wire   [0:0] icmp_ln289_fu_4792_p2;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
wire   [7:0] ap_phi_reg_pp0_iter0_act_m_val_V_reg_1636;
reg   [7:0] ap_phi_reg_pp0_iter1_act_m_val_V_reg_1636;
reg   [15:0] tmp_V_fu_570;
wire   [15:0] tmp_V_260_fu_4871_p2;
reg   [31:0] sf_1_fu_574;
wire   [31:0] sf_fu_4786_p2;
reg   [7:0] tmp_V_1_fu_578;
reg   [7:0] tmp_V_2_fu_582;
reg   [7:0] tmp_V_4_fu_586;
reg   [7:0] tmp_V_5_fu_590;
reg   [7:0] tmp_V_6_fu_594;
reg   [7:0] tmp_V_7_fu_598;
reg   [7:0] tmp_V_8_fu_602;
reg   [7:0] tmp_V_9_fu_606;
reg   [7:0] tmp_V_10_fu_610;
reg   [7:0] tmp_V_11_fu_614;
reg   [7:0] tmp_V_12_fu_618;
reg   [7:0] tmp_V_13_fu_622;
reg   [7:0] tmp_V_14_fu_626;
reg   [7:0] tmp_V_15_fu_630;
reg   [7:0] tmp_V_16_fu_634;
reg   [7:0] tmp_V_17_fu_638;
reg   [7:0] tmp_V_18_fu_642;
reg   [7:0] tmp_V_19_fu_646;
reg   [7:0] tmp_V_20_fu_650;
reg   [7:0] tmp_V_21_fu_654;
reg   [7:0] tmp_V_22_fu_658;
reg   [7:0] tmp_V_23_fu_662;
reg   [7:0] tmp_V_24_fu_666;
reg   [7:0] tmp_V_25_fu_670;
reg   [7:0] tmp_V_26_fu_674;
reg   [7:0] tmp_V_27_fu_678;
reg   [7:0] tmp_V_28_fu_682;
reg   [7:0] tmp_V_29_fu_686;
reg   [7:0] tmp_V_30_fu_690;
reg   [7:0] tmp_V_31_fu_694;
reg   [7:0] tmp_V_32_fu_698;
reg   [7:0] tmp_V_33_fu_702;
reg   [7:0] tmp_V_34_fu_706;
reg   [7:0] tmp_V_35_fu_710;
reg   [7:0] tmp_V_36_fu_714;
reg   [7:0] tmp_V_37_fu_718;
reg   [7:0] tmp_V_38_fu_722;
reg   [7:0] tmp_V_39_fu_726;
reg   [7:0] tmp_V_40_fu_730;
reg   [7:0] tmp_V_41_fu_734;
reg   [7:0] tmp_V_42_fu_738;
reg   [7:0] tmp_V_43_fu_742;
reg   [7:0] tmp_V_44_fu_746;
reg   [7:0] tmp_V_45_fu_750;
reg   [7:0] tmp_V_46_fu_754;
reg   [7:0] tmp_V_47_fu_758;
reg   [7:0] tmp_V_48_fu_762;
reg   [7:0] tmp_V_49_fu_766;
reg   [7:0] tmp_V_50_fu_770;
reg   [7:0] tmp_V_51_fu_774;
reg   [7:0] tmp_V_52_fu_778;
reg   [7:0] tmp_V_53_fu_782;
reg   [7:0] tmp_V_54_fu_786;
reg   [7:0] tmp_V_55_fu_790;
reg   [7:0] tmp_V_56_fu_794;
reg   [7:0] tmp_V_57_fu_798;
reg   [7:0] tmp_V_58_fu_802;
reg   [7:0] tmp_V_59_fu_806;
reg   [7:0] tmp_V_60_fu_810;
reg   [7:0] tmp_V_61_fu_814;
reg   [7:0] tmp_V_62_fu_818;
reg   [7:0] tmp_V_63_fu_822;
reg   [7:0] tmp_V_64_fu_826;
reg   [7:0] tmp_V_65_fu_830;
reg   [7:0] tmp_V_66_fu_834;
reg   [7:0] tmp_V_67_fu_838;
reg   [7:0] tmp_V_68_fu_842;
reg   [7:0] tmp_V_69_fu_846;
reg   [7:0] tmp_V_70_fu_850;
reg   [7:0] tmp_V_71_fu_854;
reg   [7:0] tmp_V_72_fu_858;
reg   [7:0] tmp_V_73_fu_862;
reg   [7:0] tmp_V_74_fu_866;
reg   [7:0] tmp_V_75_fu_870;
reg   [7:0] tmp_V_76_fu_874;
reg   [7:0] tmp_V_77_fu_878;
reg   [7:0] tmp_V_78_fu_882;
reg   [7:0] tmp_V_79_fu_886;
reg   [7:0] tmp_V_80_fu_890;
reg   [7:0] tmp_V_81_fu_894;
reg   [7:0] tmp_V_82_fu_898;
reg   [7:0] tmp_V_83_fu_902;
reg   [7:0] tmp_V_84_fu_906;
reg   [7:0] tmp_V_85_fu_910;
reg   [7:0] tmp_V_86_fu_914;
reg   [7:0] tmp_V_87_fu_918;
reg   [7:0] tmp_V_88_fu_922;
reg   [7:0] tmp_V_89_fu_926;
reg   [7:0] tmp_V_90_fu_930;
reg   [7:0] tmp_V_91_fu_934;
reg   [7:0] tmp_V_92_fu_938;
reg   [7:0] tmp_V_93_fu_942;
reg   [7:0] tmp_V_94_fu_946;
reg   [7:0] tmp_V_95_fu_950;
reg   [7:0] tmp_V_96_fu_954;
reg   [7:0] tmp_V_97_fu_958;
reg   [7:0] tmp_V_98_fu_962;
reg   [7:0] tmp_V_99_fu_966;
reg   [7:0] tmp_V_100_fu_970;
reg   [7:0] tmp_V_101_fu_974;
reg   [7:0] tmp_V_102_fu_978;
reg   [7:0] tmp_V_103_fu_982;
reg   [7:0] tmp_V_104_fu_986;
reg   [7:0] tmp_V_105_fu_990;
reg   [7:0] tmp_V_106_fu_994;
reg   [7:0] tmp_V_107_fu_998;
reg   [7:0] tmp_V_108_fu_1002;
reg   [7:0] tmp_V_109_fu_1006;
reg   [7:0] tmp_V_110_fu_1010;
reg   [7:0] tmp_V_111_fu_1014;
reg   [7:0] tmp_V_112_fu_1018;
reg   [7:0] tmp_V_113_fu_1022;
reg   [7:0] tmp_V_114_fu_1026;
reg   [7:0] tmp_V_115_fu_1030;
reg   [7:0] tmp_V_116_fu_1034;
reg   [7:0] tmp_V_117_fu_1038;
reg   [7:0] tmp_V_118_fu_1042;
reg   [7:0] tmp_V_119_fu_1046;
reg   [7:0] tmp_V_120_fu_1050;
reg   [7:0] tmp_V_121_fu_1054;
reg   [7:0] tmp_V_122_fu_1058;
reg   [7:0] tmp_V_123_fu_1062;
reg   [7:0] tmp_V_124_fu_1066;
reg   [7:0] tmp_V_125_fu_1070;
reg   [7:0] tmp_V_126_fu_1074;
reg   [7:0] tmp_V_127_fu_1078;
reg   [7:0] tmp_V_128_fu_1082;
reg   [7:0] tmp_V_129_fu_1086;
reg   [7:0] tmp_V_130_fu_1090;
reg   [7:0] tmp_V_131_fu_1094;
reg   [7:0] tmp_V_132_fu_1098;
reg   [7:0] tmp_V_133_fu_1102;
reg   [7:0] tmp_V_134_fu_1106;
reg   [7:0] tmp_V_135_fu_1110;
reg   [7:0] tmp_V_136_fu_1114;
reg   [7:0] tmp_V_137_fu_1118;
reg   [7:0] tmp_V_138_fu_1122;
reg   [7:0] tmp_V_139_fu_1126;
reg   [7:0] tmp_V_140_fu_1130;
reg   [7:0] tmp_V_141_fu_1134;
reg   [7:0] tmp_V_142_fu_1138;
reg   [7:0] tmp_V_143_fu_1142;
reg   [7:0] tmp_V_144_fu_1146;
reg   [7:0] tmp_V_145_fu_1150;
reg   [7:0] tmp_V_146_fu_1154;
reg   [7:0] tmp_V_147_fu_1158;
reg   [7:0] tmp_V_148_fu_1162;
reg   [7:0] tmp_V_149_fu_1166;
reg   [7:0] tmp_V_150_fu_1170;
reg   [7:0] tmp_V_151_fu_1174;
reg   [7:0] tmp_V_152_fu_1178;
reg   [7:0] tmp_V_153_fu_1182;
reg   [7:0] tmp_V_154_fu_1186;
reg   [7:0] tmp_V_155_fu_1190;
reg   [7:0] tmp_V_156_fu_1194;
reg   [7:0] tmp_V_157_fu_1198;
reg   [7:0] tmp_V_158_fu_1202;
reg   [7:0] tmp_V_159_fu_1206;
reg   [7:0] tmp_V_160_fu_1210;
reg   [7:0] tmp_V_161_fu_1214;
reg   [7:0] tmp_V_162_fu_1218;
reg   [7:0] tmp_V_163_fu_1222;
reg   [7:0] tmp_V_164_fu_1226;
reg   [7:0] tmp_V_165_fu_1230;
reg   [7:0] tmp_V_166_fu_1234;
reg   [7:0] tmp_V_167_fu_1238;
reg   [7:0] tmp_V_168_fu_1242;
reg   [7:0] tmp_V_169_fu_1246;
reg   [7:0] tmp_V_170_fu_1250;
reg   [7:0] tmp_V_171_fu_1254;
reg   [7:0] tmp_V_172_fu_1258;
reg   [7:0] tmp_V_173_fu_1262;
reg   [7:0] tmp_V_174_fu_1266;
reg   [7:0] tmp_V_175_fu_1270;
reg   [7:0] tmp_V_176_fu_1274;
reg   [7:0] tmp_V_177_fu_1278;
reg   [7:0] tmp_V_178_fu_1282;
reg   [7:0] tmp_V_179_fu_1286;
reg   [7:0] tmp_V_180_fu_1290;
reg   [7:0] tmp_V_181_fu_1294;
reg   [7:0] tmp_V_182_fu_1298;
reg   [7:0] tmp_V_183_fu_1302;
reg   [7:0] tmp_V_184_fu_1306;
reg   [7:0] tmp_V_185_fu_1310;
reg   [7:0] tmp_V_186_fu_1314;
reg   [7:0] tmp_V_187_fu_1318;
reg   [7:0] tmp_V_188_fu_1322;
reg   [7:0] tmp_V_189_fu_1326;
reg   [7:0] tmp_V_190_fu_1330;
reg   [7:0] tmp_V_191_fu_1334;
reg   [7:0] tmp_V_192_fu_1338;
reg   [7:0] tmp_V_193_fu_1342;
reg   [7:0] tmp_V_194_fu_1346;
reg   [7:0] tmp_V_195_fu_1350;
reg   [7:0] tmp_V_196_fu_1354;
reg   [7:0] tmp_V_197_fu_1358;
reg   [7:0] tmp_V_198_fu_1362;
reg   [7:0] tmp_V_199_fu_1366;
reg   [7:0] tmp_V_200_fu_1370;
reg   [7:0] tmp_V_201_fu_1374;
reg   [7:0] tmp_V_202_fu_1378;
reg   [7:0] tmp_V_203_fu_1382;
reg   [7:0] tmp_V_204_fu_1386;
reg   [7:0] tmp_V_205_fu_1390;
reg   [7:0] tmp_V_206_fu_1394;
reg   [7:0] tmp_V_207_fu_1398;
reg   [7:0] tmp_V_208_fu_1402;
reg   [7:0] tmp_V_209_fu_1406;
reg   [7:0] tmp_V_210_fu_1410;
reg   [7:0] tmp_V_211_fu_1414;
reg   [7:0] tmp_V_212_fu_1418;
reg   [7:0] tmp_V_213_fu_1422;
reg   [7:0] tmp_V_214_fu_1426;
reg   [7:0] tmp_V_215_fu_1430;
reg   [7:0] tmp_V_216_fu_1434;
reg   [7:0] tmp_V_217_fu_1438;
reg   [7:0] tmp_V_218_fu_1442;
reg   [7:0] tmp_V_219_fu_1446;
reg   [7:0] tmp_V_220_fu_1450;
reg   [7:0] tmp_V_221_fu_1454;
reg   [7:0] tmp_V_222_fu_1458;
reg   [7:0] tmp_V_223_fu_1462;
reg   [7:0] tmp_V_224_fu_1466;
reg   [7:0] tmp_V_225_fu_1470;
reg   [7:0] tmp_V_226_fu_1474;
reg   [7:0] tmp_V_227_fu_1478;
reg   [7:0] tmp_V_228_fu_1482;
reg   [7:0] tmp_V_229_fu_1486;
reg   [7:0] tmp_V_230_fu_1490;
reg   [7:0] tmp_V_231_fu_1494;
reg   [7:0] tmp_V_232_fu_1498;
reg   [7:0] tmp_V_233_fu_1502;
reg   [7:0] tmp_V_234_fu_1506;
reg   [7:0] tmp_V_235_fu_1510;
reg   [7:0] tmp_V_236_fu_1514;
reg   [7:0] tmp_V_237_fu_1518;
reg   [7:0] tmp_V_238_fu_1522;
reg   [7:0] tmp_V_239_fu_1526;
reg   [7:0] tmp_V_240_fu_1530;
reg   [7:0] tmp_V_241_fu_1534;
reg   [7:0] tmp_V_242_fu_1538;
reg   [7:0] tmp_V_243_fu_1542;
reg   [7:0] tmp_V_244_fu_1546;
reg   [7:0] tmp_V_245_fu_1550;
reg   [7:0] tmp_V_246_fu_1554;
reg   [7:0] tmp_V_247_fu_1558;
reg   [7:0] tmp_V_248_fu_1562;
reg   [7:0] tmp_V_249_fu_1566;
reg   [7:0] tmp_V_250_fu_1570;
reg   [7:0] tmp_V_251_fu_1574;
reg   [7:0] tmp_V_252_fu_1578;
reg   [7:0] tmp_V_253_fu_1582;
reg   [7:0] tmp_V_254_fu_1586;
reg   [7:0] tmp_V_255_fu_1590;
reg   [7:0] tmp_V_256_fu_1594;
reg   [7:0] tmp_V_257_fu_1598;
reg   [31:0] nf_2_fu_1602;
wire   [31:0] nf_3_fu_4898_p3;
reg   [31:0] ap_sig_allocacmp_nf_2_load;
reg    ap_block_pp0_stage0_01001;
wire   [7:0] inElem_V_1_fu_2961_p257;
wire  signed [3:0] trunc_ln647_1_fu_4813_p1;
wire  signed [7:0] mul_ln1352_fu_4824_p2;
wire  signed [3:0] arg_V_read_assign_1_fu_4834_p4;
wire  signed [7:0] mul_ln1352_1_fu_4851_p2;
wire  signed [8:0] sext_ln700_fu_4857_p1;
wire  signed [8:0] sext_ln170_fu_4830_p1;
wire   [8:0] add_ln700_fu_4861_p2;
wire   [15:0] res_V_fu_4806_p3;
wire  signed [15:0] sext_ln700_1_fu_4867_p1;
wire   [31:0] nf_fu_4886_p2;
wire   [0:0] icmp_ln301_fu_4892_p2;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

StreamingFCLayer_Batch_6_StreamingFCLayer_bkb #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 8 ),
    .din2_WIDTH( 8 ),
    .din3_WIDTH( 8 ),
    .din4_WIDTH( 8 ),
    .din5_WIDTH( 8 ),
    .din6_WIDTH( 8 ),
    .din7_WIDTH( 8 ),
    .din8_WIDTH( 8 ),
    .din9_WIDTH( 8 ),
    .din10_WIDTH( 8 ),
    .din11_WIDTH( 8 ),
    .din12_WIDTH( 8 ),
    .din13_WIDTH( 8 ),
    .din14_WIDTH( 8 ),
    .din15_WIDTH( 8 ),
    .din16_WIDTH( 8 ),
    .din17_WIDTH( 8 ),
    .din18_WIDTH( 8 ),
    .din19_WIDTH( 8 ),
    .din20_WIDTH( 8 ),
    .din21_WIDTH( 8 ),
    .din22_WIDTH( 8 ),
    .din23_WIDTH( 8 ),
    .din24_WIDTH( 8 ),
    .din25_WIDTH( 8 ),
    .din26_WIDTH( 8 ),
    .din27_WIDTH( 8 ),
    .din28_WIDTH( 8 ),
    .din29_WIDTH( 8 ),
    .din30_WIDTH( 8 ),
    .din31_WIDTH( 8 ),
    .din32_WIDTH( 8 ),
    .din33_WIDTH( 8 ),
    .din34_WIDTH( 8 ),
    .din35_WIDTH( 8 ),
    .din36_WIDTH( 8 ),
    .din37_WIDTH( 8 ),
    .din38_WIDTH( 8 ),
    .din39_WIDTH( 8 ),
    .din40_WIDTH( 8 ),
    .din41_WIDTH( 8 ),
    .din42_WIDTH( 8 ),
    .din43_WIDTH( 8 ),
    .din44_WIDTH( 8 ),
    .din45_WIDTH( 8 ),
    .din46_WIDTH( 8 ),
    .din47_WIDTH( 8 ),
    .din48_WIDTH( 8 ),
    .din49_WIDTH( 8 ),
    .din50_WIDTH( 8 ),
    .din51_WIDTH( 8 ),
    .din52_WIDTH( 8 ),
    .din53_WIDTH( 8 ),
    .din54_WIDTH( 8 ),
    .din55_WIDTH( 8 ),
    .din56_WIDTH( 8 ),
    .din57_WIDTH( 8 ),
    .din58_WIDTH( 8 ),
    .din59_WIDTH( 8 ),
    .din60_WIDTH( 8 ),
    .din61_WIDTH( 8 ),
    .din62_WIDTH( 8 ),
    .din63_WIDTH( 8 ),
    .din64_WIDTH( 8 ),
    .din65_WIDTH( 8 ),
    .din66_WIDTH( 8 ),
    .din67_WIDTH( 8 ),
    .din68_WIDTH( 8 ),
    .din69_WIDTH( 8 ),
    .din70_WIDTH( 8 ),
    .din71_WIDTH( 8 ),
    .din72_WIDTH( 8 ),
    .din73_WIDTH( 8 ),
    .din74_WIDTH( 8 ),
    .din75_WIDTH( 8 ),
    .din76_WIDTH( 8 ),
    .din77_WIDTH( 8 ),
    .din78_WIDTH( 8 ),
    .din79_WIDTH( 8 ),
    .din80_WIDTH( 8 ),
    .din81_WIDTH( 8 ),
    .din82_WIDTH( 8 ),
    .din83_WIDTH( 8 ),
    .din84_WIDTH( 8 ),
    .din85_WIDTH( 8 ),
    .din86_WIDTH( 8 ),
    .din87_WIDTH( 8 ),
    .din88_WIDTH( 8 ),
    .din89_WIDTH( 8 ),
    .din90_WIDTH( 8 ),
    .din91_WIDTH( 8 ),
    .din92_WIDTH( 8 ),
    .din93_WIDTH( 8 ),
    .din94_WIDTH( 8 ),
    .din95_WIDTH( 8 ),
    .din96_WIDTH( 8 ),
    .din97_WIDTH( 8 ),
    .din98_WIDTH( 8 ),
    .din99_WIDTH( 8 ),
    .din100_WIDTH( 8 ),
    .din101_WIDTH( 8 ),
    .din102_WIDTH( 8 ),
    .din103_WIDTH( 8 ),
    .din104_WIDTH( 8 ),
    .din105_WIDTH( 8 ),
    .din106_WIDTH( 8 ),
    .din107_WIDTH( 8 ),
    .din108_WIDTH( 8 ),
    .din109_WIDTH( 8 ),
    .din110_WIDTH( 8 ),
    .din111_WIDTH( 8 ),
    .din112_WIDTH( 8 ),
    .din113_WIDTH( 8 ),
    .din114_WIDTH( 8 ),
    .din115_WIDTH( 8 ),
    .din116_WIDTH( 8 ),
    .din117_WIDTH( 8 ),
    .din118_WIDTH( 8 ),
    .din119_WIDTH( 8 ),
    .din120_WIDTH( 8 ),
    .din121_WIDTH( 8 ),
    .din122_WIDTH( 8 ),
    .din123_WIDTH( 8 ),
    .din124_WIDTH( 8 ),
    .din125_WIDTH( 8 ),
    .din126_WIDTH( 8 ),
    .din127_WIDTH( 8 ),
    .din128_WIDTH( 8 ),
    .din129_WIDTH( 8 ),
    .din130_WIDTH( 8 ),
    .din131_WIDTH( 8 ),
    .din132_WIDTH( 8 ),
    .din133_WIDTH( 8 ),
    .din134_WIDTH( 8 ),
    .din135_WIDTH( 8 ),
    .din136_WIDTH( 8 ),
    .din137_WIDTH( 8 ),
    .din138_WIDTH( 8 ),
    .din139_WIDTH( 8 ),
    .din140_WIDTH( 8 ),
    .din141_WIDTH( 8 ),
    .din142_WIDTH( 8 ),
    .din143_WIDTH( 8 ),
    .din144_WIDTH( 8 ),
    .din145_WIDTH( 8 ),
    .din146_WIDTH( 8 ),
    .din147_WIDTH( 8 ),
    .din148_WIDTH( 8 ),
    .din149_WIDTH( 8 ),
    .din150_WIDTH( 8 ),
    .din151_WIDTH( 8 ),
    .din152_WIDTH( 8 ),
    .din153_WIDTH( 8 ),
    .din154_WIDTH( 8 ),
    .din155_WIDTH( 8 ),
    .din156_WIDTH( 8 ),
    .din157_WIDTH( 8 ),
    .din158_WIDTH( 8 ),
    .din159_WIDTH( 8 ),
    .din160_WIDTH( 8 ),
    .din161_WIDTH( 8 ),
    .din162_WIDTH( 8 ),
    .din163_WIDTH( 8 ),
    .din164_WIDTH( 8 ),
    .din165_WIDTH( 8 ),
    .din166_WIDTH( 8 ),
    .din167_WIDTH( 8 ),
    .din168_WIDTH( 8 ),
    .din169_WIDTH( 8 ),
    .din170_WIDTH( 8 ),
    .din171_WIDTH( 8 ),
    .din172_WIDTH( 8 ),
    .din173_WIDTH( 8 ),
    .din174_WIDTH( 8 ),
    .din175_WIDTH( 8 ),
    .din176_WIDTH( 8 ),
    .din177_WIDTH( 8 ),
    .din178_WIDTH( 8 ),
    .din179_WIDTH( 8 ),
    .din180_WIDTH( 8 ),
    .din181_WIDTH( 8 ),
    .din182_WIDTH( 8 ),
    .din183_WIDTH( 8 ),
    .din184_WIDTH( 8 ),
    .din185_WIDTH( 8 ),
    .din186_WIDTH( 8 ),
    .din187_WIDTH( 8 ),
    .din188_WIDTH( 8 ),
    .din189_WIDTH( 8 ),
    .din190_WIDTH( 8 ),
    .din191_WIDTH( 8 ),
    .din192_WIDTH( 8 ),
    .din193_WIDTH( 8 ),
    .din194_WIDTH( 8 ),
    .din195_WIDTH( 8 ),
    .din196_WIDTH( 8 ),
    .din197_WIDTH( 8 ),
    .din198_WIDTH( 8 ),
    .din199_WIDTH( 8 ),
    .din200_WIDTH( 8 ),
    .din201_WIDTH( 8 ),
    .din202_WIDTH( 8 ),
    .din203_WIDTH( 8 ),
    .din204_WIDTH( 8 ),
    .din205_WIDTH( 8 ),
    .din206_WIDTH( 8 ),
    .din207_WIDTH( 8 ),
    .din208_WIDTH( 8 ),
    .din209_WIDTH( 8 ),
    .din210_WIDTH( 8 ),
    .din211_WIDTH( 8 ),
    .din212_WIDTH( 8 ),
    .din213_WIDTH( 8 ),
    .din214_WIDTH( 8 ),
    .din215_WIDTH( 8 ),
    .din216_WIDTH( 8 ),
    .din217_WIDTH( 8 ),
    .din218_WIDTH( 8 ),
    .din219_WIDTH( 8 ),
    .din220_WIDTH( 8 ),
    .din221_WIDTH( 8 ),
    .din222_WIDTH( 8 ),
    .din223_WIDTH( 8 ),
    .din224_WIDTH( 8 ),
    .din225_WIDTH( 8 ),
    .din226_WIDTH( 8 ),
    .din227_WIDTH( 8 ),
    .din228_WIDTH( 8 ),
    .din229_WIDTH( 8 ),
    .din230_WIDTH( 8 ),
    .din231_WIDTH( 8 ),
    .din232_WIDTH( 8 ),
    .din233_WIDTH( 8 ),
    .din234_WIDTH( 8 ),
    .din235_WIDTH( 8 ),
    .din236_WIDTH( 8 ),
    .din237_WIDTH( 8 ),
    .din238_WIDTH( 8 ),
    .din239_WIDTH( 8 ),
    .din240_WIDTH( 8 ),
    .din241_WIDTH( 8 ),
    .din242_WIDTH( 8 ),
    .din243_WIDTH( 8 ),
    .din244_WIDTH( 8 ),
    .din245_WIDTH( 8 ),
    .din246_WIDTH( 8 ),
    .din247_WIDTH( 8 ),
    .din248_WIDTH( 8 ),
    .din249_WIDTH( 8 ),
    .din250_WIDTH( 8 ),
    .din251_WIDTH( 8 ),
    .din252_WIDTH( 8 ),
    .din253_WIDTH( 8 ),
    .din254_WIDTH( 8 ),
    .din255_WIDTH( 8 ),
    .din256_WIDTH( 8 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_bkb_U1(
    .din0(tmp_V_1_fu_578),
    .din1(tmp_V_2_fu_582),
    .din2(tmp_V_4_fu_586),
    .din3(tmp_V_5_fu_590),
    .din4(tmp_V_6_fu_594),
    .din5(tmp_V_7_fu_598),
    .din6(tmp_V_8_fu_602),
    .din7(tmp_V_9_fu_606),
    .din8(tmp_V_10_fu_610),
    .din9(tmp_V_11_fu_614),
    .din10(tmp_V_12_fu_618),
    .din11(tmp_V_13_fu_622),
    .din12(tmp_V_14_fu_626),
    .din13(tmp_V_15_fu_630),
    .din14(tmp_V_16_fu_634),
    .din15(tmp_V_17_fu_638),
    .din16(tmp_V_18_fu_642),
    .din17(tmp_V_19_fu_646),
    .din18(tmp_V_20_fu_650),
    .din19(tmp_V_21_fu_654),
    .din20(tmp_V_22_fu_658),
    .din21(tmp_V_23_fu_662),
    .din22(tmp_V_24_fu_666),
    .din23(tmp_V_25_fu_670),
    .din24(tmp_V_26_fu_674),
    .din25(tmp_V_27_fu_678),
    .din26(tmp_V_28_fu_682),
    .din27(tmp_V_29_fu_686),
    .din28(tmp_V_30_fu_690),
    .din29(tmp_V_31_fu_694),
    .din30(tmp_V_32_fu_698),
    .din31(tmp_V_33_fu_702),
    .din32(tmp_V_34_fu_706),
    .din33(tmp_V_35_fu_710),
    .din34(tmp_V_36_fu_714),
    .din35(tmp_V_37_fu_718),
    .din36(tmp_V_38_fu_722),
    .din37(tmp_V_39_fu_726),
    .din38(tmp_V_40_fu_730),
    .din39(tmp_V_41_fu_734),
    .din40(tmp_V_42_fu_738),
    .din41(tmp_V_43_fu_742),
    .din42(tmp_V_44_fu_746),
    .din43(tmp_V_45_fu_750),
    .din44(tmp_V_46_fu_754),
    .din45(tmp_V_47_fu_758),
    .din46(tmp_V_48_fu_762),
    .din47(tmp_V_49_fu_766),
    .din48(tmp_V_50_fu_770),
    .din49(tmp_V_51_fu_774),
    .din50(tmp_V_52_fu_778),
    .din51(tmp_V_53_fu_782),
    .din52(tmp_V_54_fu_786),
    .din53(tmp_V_55_fu_790),
    .din54(tmp_V_56_fu_794),
    .din55(tmp_V_57_fu_798),
    .din56(tmp_V_58_fu_802),
    .din57(tmp_V_59_fu_806),
    .din58(tmp_V_60_fu_810),
    .din59(tmp_V_61_fu_814),
    .din60(tmp_V_62_fu_818),
    .din61(tmp_V_63_fu_822),
    .din62(tmp_V_64_fu_826),
    .din63(tmp_V_65_fu_830),
    .din64(tmp_V_66_fu_834),
    .din65(tmp_V_67_fu_838),
    .din66(tmp_V_68_fu_842),
    .din67(tmp_V_69_fu_846),
    .din68(tmp_V_70_fu_850),
    .din69(tmp_V_71_fu_854),
    .din70(tmp_V_72_fu_858),
    .din71(tmp_V_73_fu_862),
    .din72(tmp_V_74_fu_866),
    .din73(tmp_V_75_fu_870),
    .din74(tmp_V_76_fu_874),
    .din75(tmp_V_77_fu_878),
    .din76(tmp_V_78_fu_882),
    .din77(tmp_V_79_fu_886),
    .din78(tmp_V_80_fu_890),
    .din79(tmp_V_81_fu_894),
    .din80(tmp_V_82_fu_898),
    .din81(tmp_V_83_fu_902),
    .din82(tmp_V_84_fu_906),
    .din83(tmp_V_85_fu_910),
    .din84(tmp_V_86_fu_914),
    .din85(tmp_V_87_fu_918),
    .din86(tmp_V_88_fu_922),
    .din87(tmp_V_89_fu_926),
    .din88(tmp_V_90_fu_930),
    .din89(tmp_V_91_fu_934),
    .din90(tmp_V_92_fu_938),
    .din91(tmp_V_93_fu_942),
    .din92(tmp_V_94_fu_946),
    .din93(tmp_V_95_fu_950),
    .din94(tmp_V_96_fu_954),
    .din95(tmp_V_97_fu_958),
    .din96(tmp_V_98_fu_962),
    .din97(tmp_V_99_fu_966),
    .din98(tmp_V_100_fu_970),
    .din99(tmp_V_101_fu_974),
    .din100(tmp_V_102_fu_978),
    .din101(tmp_V_103_fu_982),
    .din102(tmp_V_104_fu_986),
    .din103(tmp_V_105_fu_990),
    .din104(tmp_V_106_fu_994),
    .din105(tmp_V_107_fu_998),
    .din106(tmp_V_108_fu_1002),
    .din107(tmp_V_109_fu_1006),
    .din108(tmp_V_110_fu_1010),
    .din109(tmp_V_111_fu_1014),
    .din110(tmp_V_112_fu_1018),
    .din111(tmp_V_113_fu_1022),
    .din112(tmp_V_114_fu_1026),
    .din113(tmp_V_115_fu_1030),
    .din114(tmp_V_116_fu_1034),
    .din115(tmp_V_117_fu_1038),
    .din116(tmp_V_118_fu_1042),
    .din117(tmp_V_119_fu_1046),
    .din118(tmp_V_120_fu_1050),
    .din119(tmp_V_121_fu_1054),
    .din120(tmp_V_122_fu_1058),
    .din121(tmp_V_123_fu_1062),
    .din122(tmp_V_124_fu_1066),
    .din123(tmp_V_125_fu_1070),
    .din124(tmp_V_126_fu_1074),
    .din125(tmp_V_127_fu_1078),
    .din126(tmp_V_128_fu_1082),
    .din127(tmp_V_129_fu_1086),
    .din128(tmp_V_130_fu_1090),
    .din129(tmp_V_131_fu_1094),
    .din130(tmp_V_132_fu_1098),
    .din131(tmp_V_133_fu_1102),
    .din132(tmp_V_134_fu_1106),
    .din133(tmp_V_135_fu_1110),
    .din134(tmp_V_136_fu_1114),
    .din135(tmp_V_137_fu_1118),
    .din136(tmp_V_138_fu_1122),
    .din137(tmp_V_139_fu_1126),
    .din138(tmp_V_140_fu_1130),
    .din139(tmp_V_141_fu_1134),
    .din140(tmp_V_142_fu_1138),
    .din141(tmp_V_143_fu_1142),
    .din142(tmp_V_144_fu_1146),
    .din143(tmp_V_145_fu_1150),
    .din144(tmp_V_146_fu_1154),
    .din145(tmp_V_147_fu_1158),
    .din146(tmp_V_148_fu_1162),
    .din147(tmp_V_149_fu_1166),
    .din148(tmp_V_150_fu_1170),
    .din149(tmp_V_151_fu_1174),
    .din150(tmp_V_152_fu_1178),
    .din151(tmp_V_153_fu_1182),
    .din152(tmp_V_154_fu_1186),
    .din153(tmp_V_155_fu_1190),
    .din154(tmp_V_156_fu_1194),
    .din155(tmp_V_157_fu_1198),
    .din156(tmp_V_158_fu_1202),
    .din157(tmp_V_159_fu_1206),
    .din158(tmp_V_160_fu_1210),
    .din159(tmp_V_161_fu_1214),
    .din160(tmp_V_162_fu_1218),
    .din161(tmp_V_163_fu_1222),
    .din162(tmp_V_164_fu_1226),
    .din163(tmp_V_165_fu_1230),
    .din164(tmp_V_166_fu_1234),
    .din165(tmp_V_167_fu_1238),
    .din166(tmp_V_168_fu_1242),
    .din167(tmp_V_169_fu_1246),
    .din168(tmp_V_170_fu_1250),
    .din169(tmp_V_171_fu_1254),
    .din170(tmp_V_172_fu_1258),
    .din171(tmp_V_173_fu_1262),
    .din172(tmp_V_174_fu_1266),
    .din173(tmp_V_175_fu_1270),
    .din174(tmp_V_176_fu_1274),
    .din175(tmp_V_177_fu_1278),
    .din176(tmp_V_178_fu_1282),
    .din177(tmp_V_179_fu_1286),
    .din178(tmp_V_180_fu_1290),
    .din179(tmp_V_181_fu_1294),
    .din180(tmp_V_182_fu_1298),
    .din181(tmp_V_183_fu_1302),
    .din182(tmp_V_184_fu_1306),
    .din183(tmp_V_185_fu_1310),
    .din184(tmp_V_186_fu_1314),
    .din185(tmp_V_187_fu_1318),
    .din186(tmp_V_188_fu_1322),
    .din187(tmp_V_189_fu_1326),
    .din188(tmp_V_190_fu_1330),
    .din189(tmp_V_191_fu_1334),
    .din190(tmp_V_192_fu_1338),
    .din191(tmp_V_193_fu_1342),
    .din192(tmp_V_194_fu_1346),
    .din193(tmp_V_195_fu_1350),
    .din194(tmp_V_196_fu_1354),
    .din195(tmp_V_197_fu_1358),
    .din196(tmp_V_198_fu_1362),
    .din197(tmp_V_199_fu_1366),
    .din198(tmp_V_200_fu_1370),
    .din199(tmp_V_201_fu_1374),
    .din200(tmp_V_202_fu_1378),
    .din201(tmp_V_203_fu_1382),
    .din202(tmp_V_204_fu_1386),
    .din203(tmp_V_205_fu_1390),
    .din204(tmp_V_206_fu_1394),
    .din205(tmp_V_207_fu_1398),
    .din206(tmp_V_208_fu_1402),
    .din207(tmp_V_209_fu_1406),
    .din208(tmp_V_210_fu_1410),
    .din209(tmp_V_211_fu_1414),
    .din210(tmp_V_212_fu_1418),
    .din211(tmp_V_213_fu_1422),
    .din212(tmp_V_214_fu_1426),
    .din213(tmp_V_215_fu_1430),
    .din214(tmp_V_216_fu_1434),
    .din215(tmp_V_217_fu_1438),
    .din216(tmp_V_218_fu_1442),
    .din217(tmp_V_219_fu_1446),
    .din218(tmp_V_220_fu_1450),
    .din219(tmp_V_221_fu_1454),
    .din220(tmp_V_222_fu_1458),
    .din221(tmp_V_223_fu_1462),
    .din222(tmp_V_224_fu_1466),
    .din223(tmp_V_225_fu_1470),
    .din224(tmp_V_226_fu_1474),
    .din225(tmp_V_227_fu_1478),
    .din226(tmp_V_228_fu_1482),
    .din227(tmp_V_229_fu_1486),
    .din228(tmp_V_230_fu_1490),
    .din229(tmp_V_231_fu_1494),
    .din230(tmp_V_232_fu_1498),
    .din231(tmp_V_233_fu_1502),
    .din232(tmp_V_234_fu_1506),
    .din233(tmp_V_235_fu_1510),
    .din234(tmp_V_236_fu_1514),
    .din235(tmp_V_237_fu_1518),
    .din236(tmp_V_238_fu_1522),
    .din237(tmp_V_239_fu_1526),
    .din238(tmp_V_240_fu_1530),
    .din239(tmp_V_241_fu_1534),
    .din240(tmp_V_242_fu_1538),
    .din241(tmp_V_243_fu_1542),
    .din242(tmp_V_244_fu_1546),
    .din243(tmp_V_245_fu_1550),
    .din244(tmp_V_246_fu_1554),
    .din245(tmp_V_247_fu_1558),
    .din246(tmp_V_248_fu_1562),
    .din247(tmp_V_249_fu_1566),
    .din248(tmp_V_250_fu_1570),
    .din249(tmp_V_251_fu_1574),
    .din250(tmp_V_252_fu_1578),
    .din251(tmp_V_253_fu_1582),
    .din252(tmp_V_254_fu_1586),
    .din253(tmp_V_255_fu_1590),
    .din254(tmp_V_256_fu_1594),
    .din255(tmp_V_257_fu_1598),
    .din256(inElem_V_1_fu_2961_p257),
    .dout(inElem_V_1_fu_2961_p258)
);

StreamingFCLayer_Batch_6_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U2(
    .din0(trunc_ln647_1_fu_4813_p1),
    .din1(trunc_ln647_reg_6756),
    .dout(mul_ln1352_fu_4824_p2)
);

StreamingFCLayer_Batch_6_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U3(
    .din0(arg_V_read_assign_1_fu_4834_p4),
    .din1(p_Result_s_reg_6761),
    .dout(mul_ln1352_1_fu_4851_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd0) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_1636 <= inElem_V_1_fu_2961_p258;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd82)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd83)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd84)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd85)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd86)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd87)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd88)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd89)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd90)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd91)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd92)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd93)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd94)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd95)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd96)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd97)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd98)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd99)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd100)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd101)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd102)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd103)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd104)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd105)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd106)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd107)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd108)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd109)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd110)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd111)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd112)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd113)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd114)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd115)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd116)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd117)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd118)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd119)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd120)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd121)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd122)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd123)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd124)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd125)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd126)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd127)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd128)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd129)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd130)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd131)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd132)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd133)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd134)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd135)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd136)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd137)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd138)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd139)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd140)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd141)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd142)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd143)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd144)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd145)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd146)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd147)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd148)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd149)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd150)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd151)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd152)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd153)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd154)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd155)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd156)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd157)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd158)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd159)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd160)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd161)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd162)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd163)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd164)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd165)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd166)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd167)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd168)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd169)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd170)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd171)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd172)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd173)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd174)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd175)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd176)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd177)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd178)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd179)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd180)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd181)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd182)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd183)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd184)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd185)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd186)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd187)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd188)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd189)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd190)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd191)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd192)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd193)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd194)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd195)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd196)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd197)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd198)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd199)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd200)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd201)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd202)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd203)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd204)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd205)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd206)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd207)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd208)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd209)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd210)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd211)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd212)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd213)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd214)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd215)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd216)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd217)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd218)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd219)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd220)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd221)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd222)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd223)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd224)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd225)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd226)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd227)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd228)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd229)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd230)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd231)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd232)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd233)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd234)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd235)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd236)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd237)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd238)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd239)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd240)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd241)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd242)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd243)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd244)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd245)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd246)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd247)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd248)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd249)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd250)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd251)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd252)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd253)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd2)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd3)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd4)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd5)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd6)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd7)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd8)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd9)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd254)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd10)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd11)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd12)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd13)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd14)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd15)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd16)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd17)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd18)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd19)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd255)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd20)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd21)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd22)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd23)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd24)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd25)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd26)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd27)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd28)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd29)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd30)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd31)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd32)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd33)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd34)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd35)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd36)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd37)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd38)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd39)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd40)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd41)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd42)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd43)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd44)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd45)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd46)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd47)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd48)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd49)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd50)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd51)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd52)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd53)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd54)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd55)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd56)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd57)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd58)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd59)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd60)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd61)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd62)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd63)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd64)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd65)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd66)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd67)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd68)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd69)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd70)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd71)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd72)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd73)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd74)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd75)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd76)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd77)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd78)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd79)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd80)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd81)))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_1636 <= in_V_V_TDATA;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_1636 <= ap_phi_reg_pp0_iter0_act_m_val_V_reg_1636;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_reg_1625 <= i_fu_2171_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_reg_1625 <= 11'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_6766 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        nf_2_fu_1602 <= nf_3_fu_4898_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        nf_2_fu_1602 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_4792_p2 == 1'd0) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        sf_1_fu_574 <= sf_fu_4786_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_4792_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        sf_1_fu_574 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_2165_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln271_reg_6751 <= icmp_ln271_fu_4766_p2;
        icmp_ln289_reg_6766 <= icmp_ln289_fu_4792_p2;
        p_Result_s_reg_6761 <= {{weight_V_V_TDATA[7:4]}};
        trunc_ln647_reg_6756 <= trunc_ln647_fu_4772_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd98))) begin
        tmp_V_100_fu_970 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd99))) begin
        tmp_V_101_fu_974 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd100))) begin
        tmp_V_102_fu_978 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd101))) begin
        tmp_V_103_fu_982 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd102))) begin
        tmp_V_104_fu_986 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd103))) begin
        tmp_V_105_fu_990 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd104))) begin
        tmp_V_106_fu_994 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd105))) begin
        tmp_V_107_fu_998 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd106))) begin
        tmp_V_108_fu_1002 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd107))) begin
        tmp_V_109_fu_1006 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd8))) begin
        tmp_V_10_fu_610 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd108))) begin
        tmp_V_110_fu_1010 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd109))) begin
        tmp_V_111_fu_1014 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd110))) begin
        tmp_V_112_fu_1018 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd111))) begin
        tmp_V_113_fu_1022 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd112))) begin
        tmp_V_114_fu_1026 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd113))) begin
        tmp_V_115_fu_1030 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd114))) begin
        tmp_V_116_fu_1034 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd115))) begin
        tmp_V_117_fu_1038 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd116))) begin
        tmp_V_118_fu_1042 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd117))) begin
        tmp_V_119_fu_1046 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd9))) begin
        tmp_V_11_fu_614 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd118))) begin
        tmp_V_120_fu_1050 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd119))) begin
        tmp_V_121_fu_1054 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd120))) begin
        tmp_V_122_fu_1058 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd121))) begin
        tmp_V_123_fu_1062 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd122))) begin
        tmp_V_124_fu_1066 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd123))) begin
        tmp_V_125_fu_1070 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd124))) begin
        tmp_V_126_fu_1074 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd125))) begin
        tmp_V_127_fu_1078 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd126))) begin
        tmp_V_128_fu_1082 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd127))) begin
        tmp_V_129_fu_1086 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd10))) begin
        tmp_V_12_fu_618 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd128))) begin
        tmp_V_130_fu_1090 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd129))) begin
        tmp_V_131_fu_1094 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd130))) begin
        tmp_V_132_fu_1098 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd131))) begin
        tmp_V_133_fu_1102 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd132))) begin
        tmp_V_134_fu_1106 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd133))) begin
        tmp_V_135_fu_1110 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd134))) begin
        tmp_V_136_fu_1114 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd135))) begin
        tmp_V_137_fu_1118 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd136))) begin
        tmp_V_138_fu_1122 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd137))) begin
        tmp_V_139_fu_1126 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd11))) begin
        tmp_V_13_fu_622 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd138))) begin
        tmp_V_140_fu_1130 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd139))) begin
        tmp_V_141_fu_1134 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd140))) begin
        tmp_V_142_fu_1138 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd141))) begin
        tmp_V_143_fu_1142 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd142))) begin
        tmp_V_144_fu_1146 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd143))) begin
        tmp_V_145_fu_1150 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd144))) begin
        tmp_V_146_fu_1154 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd145))) begin
        tmp_V_147_fu_1158 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd146))) begin
        tmp_V_148_fu_1162 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd147))) begin
        tmp_V_149_fu_1166 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd12))) begin
        tmp_V_14_fu_626 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd148))) begin
        tmp_V_150_fu_1170 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd149))) begin
        tmp_V_151_fu_1174 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd150))) begin
        tmp_V_152_fu_1178 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd151))) begin
        tmp_V_153_fu_1182 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd152))) begin
        tmp_V_154_fu_1186 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd153))) begin
        tmp_V_155_fu_1190 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd154))) begin
        tmp_V_156_fu_1194 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd155))) begin
        tmp_V_157_fu_1198 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd156))) begin
        tmp_V_158_fu_1202 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd157))) begin
        tmp_V_159_fu_1206 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd13))) begin
        tmp_V_15_fu_630 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd158))) begin
        tmp_V_160_fu_1210 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd159))) begin
        tmp_V_161_fu_1214 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd160))) begin
        tmp_V_162_fu_1218 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd161))) begin
        tmp_V_163_fu_1222 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd162))) begin
        tmp_V_164_fu_1226 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd163))) begin
        tmp_V_165_fu_1230 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd164))) begin
        tmp_V_166_fu_1234 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd165))) begin
        tmp_V_167_fu_1238 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd166))) begin
        tmp_V_168_fu_1242 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd167))) begin
        tmp_V_169_fu_1246 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd14))) begin
        tmp_V_16_fu_634 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd168))) begin
        tmp_V_170_fu_1250 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd169))) begin
        tmp_V_171_fu_1254 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd170))) begin
        tmp_V_172_fu_1258 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd171))) begin
        tmp_V_173_fu_1262 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd172))) begin
        tmp_V_174_fu_1266 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd173))) begin
        tmp_V_175_fu_1270 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd174))) begin
        tmp_V_176_fu_1274 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd175))) begin
        tmp_V_177_fu_1278 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd176))) begin
        tmp_V_178_fu_1282 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd177))) begin
        tmp_V_179_fu_1286 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd15))) begin
        tmp_V_17_fu_638 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd178))) begin
        tmp_V_180_fu_1290 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd179))) begin
        tmp_V_181_fu_1294 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd180))) begin
        tmp_V_182_fu_1298 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd181))) begin
        tmp_V_183_fu_1302 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd182))) begin
        tmp_V_184_fu_1306 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd183))) begin
        tmp_V_185_fu_1310 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd184))) begin
        tmp_V_186_fu_1314 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd185))) begin
        tmp_V_187_fu_1318 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd186))) begin
        tmp_V_188_fu_1322 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd187))) begin
        tmp_V_189_fu_1326 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd16))) begin
        tmp_V_18_fu_642 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd188))) begin
        tmp_V_190_fu_1330 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd189))) begin
        tmp_V_191_fu_1334 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd190))) begin
        tmp_V_192_fu_1338 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd191))) begin
        tmp_V_193_fu_1342 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd192))) begin
        tmp_V_194_fu_1346 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd193))) begin
        tmp_V_195_fu_1350 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd194))) begin
        tmp_V_196_fu_1354 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd195))) begin
        tmp_V_197_fu_1358 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd196))) begin
        tmp_V_198_fu_1362 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd197))) begin
        tmp_V_199_fu_1366 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd17))) begin
        tmp_V_19_fu_646 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd0))) begin
        tmp_V_1_fu_578 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd198))) begin
        tmp_V_200_fu_1370 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd199))) begin
        tmp_V_201_fu_1374 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd200))) begin
        tmp_V_202_fu_1378 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd201))) begin
        tmp_V_203_fu_1382 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd202))) begin
        tmp_V_204_fu_1386 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd203))) begin
        tmp_V_205_fu_1390 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd204))) begin
        tmp_V_206_fu_1394 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd205))) begin
        tmp_V_207_fu_1398 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd206))) begin
        tmp_V_208_fu_1402 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd207))) begin
        tmp_V_209_fu_1406 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd18))) begin
        tmp_V_20_fu_650 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd208))) begin
        tmp_V_210_fu_1410 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd209))) begin
        tmp_V_211_fu_1414 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd210))) begin
        tmp_V_212_fu_1418 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd211))) begin
        tmp_V_213_fu_1422 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd212))) begin
        tmp_V_214_fu_1426 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd213))) begin
        tmp_V_215_fu_1430 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd214))) begin
        tmp_V_216_fu_1434 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd215))) begin
        tmp_V_217_fu_1438 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd216))) begin
        tmp_V_218_fu_1442 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd217))) begin
        tmp_V_219_fu_1446 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd19))) begin
        tmp_V_21_fu_654 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd218))) begin
        tmp_V_220_fu_1450 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd219))) begin
        tmp_V_221_fu_1454 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd220))) begin
        tmp_V_222_fu_1458 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd221))) begin
        tmp_V_223_fu_1462 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd222))) begin
        tmp_V_224_fu_1466 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd223))) begin
        tmp_V_225_fu_1470 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd224))) begin
        tmp_V_226_fu_1474 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd225))) begin
        tmp_V_227_fu_1478 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd226))) begin
        tmp_V_228_fu_1482 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd227))) begin
        tmp_V_229_fu_1486 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd20))) begin
        tmp_V_22_fu_658 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd228))) begin
        tmp_V_230_fu_1490 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd229))) begin
        tmp_V_231_fu_1494 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd230))) begin
        tmp_V_232_fu_1498 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd231))) begin
        tmp_V_233_fu_1502 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd232))) begin
        tmp_V_234_fu_1506 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd233))) begin
        tmp_V_235_fu_1510 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd234))) begin
        tmp_V_236_fu_1514 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd235))) begin
        tmp_V_237_fu_1518 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd236))) begin
        tmp_V_238_fu_1522 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd237))) begin
        tmp_V_239_fu_1526 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd21))) begin
        tmp_V_23_fu_662 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd238))) begin
        tmp_V_240_fu_1530 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd239))) begin
        tmp_V_241_fu_1534 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd240))) begin
        tmp_V_242_fu_1538 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd241))) begin
        tmp_V_243_fu_1542 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd242))) begin
        tmp_V_244_fu_1546 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd243))) begin
        tmp_V_245_fu_1550 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd244))) begin
        tmp_V_246_fu_1554 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd245))) begin
        tmp_V_247_fu_1558 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd246))) begin
        tmp_V_248_fu_1562 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd247))) begin
        tmp_V_249_fu_1566 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd22))) begin
        tmp_V_24_fu_666 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd248))) begin
        tmp_V_250_fu_1570 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd249))) begin
        tmp_V_251_fu_1574 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd250))) begin
        tmp_V_252_fu_1578 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd251))) begin
        tmp_V_253_fu_1582 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd252))) begin
        tmp_V_254_fu_1586 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd253))) begin
        tmp_V_255_fu_1590 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd254))) begin
        tmp_V_256_fu_1594 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd255))) begin
        tmp_V_257_fu_1598 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd23))) begin
        tmp_V_25_fu_670 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd24))) begin
        tmp_V_26_fu_674 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd25))) begin
        tmp_V_27_fu_678 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd26))) begin
        tmp_V_28_fu_682 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd27))) begin
        tmp_V_29_fu_686 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd1))) begin
        tmp_V_2_fu_582 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd28))) begin
        tmp_V_30_fu_690 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd29))) begin
        tmp_V_31_fu_694 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd30))) begin
        tmp_V_32_fu_698 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd31))) begin
        tmp_V_33_fu_702 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd32))) begin
        tmp_V_34_fu_706 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd33))) begin
        tmp_V_35_fu_710 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd34))) begin
        tmp_V_36_fu_714 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd35))) begin
        tmp_V_37_fu_718 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd36))) begin
        tmp_V_38_fu_722 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd37))) begin
        tmp_V_39_fu_726 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd38))) begin
        tmp_V_40_fu_730 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd39))) begin
        tmp_V_41_fu_734 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd40))) begin
        tmp_V_42_fu_738 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd41))) begin
        tmp_V_43_fu_742 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd42))) begin
        tmp_V_44_fu_746 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd43))) begin
        tmp_V_45_fu_750 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd44))) begin
        tmp_V_46_fu_754 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd45))) begin
        tmp_V_47_fu_758 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd46))) begin
        tmp_V_48_fu_762 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd47))) begin
        tmp_V_49_fu_766 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd2))) begin
        tmp_V_4_fu_586 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd48))) begin
        tmp_V_50_fu_770 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd49))) begin
        tmp_V_51_fu_774 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd50))) begin
        tmp_V_52_fu_778 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd51))) begin
        tmp_V_53_fu_782 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd52))) begin
        tmp_V_54_fu_786 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd53))) begin
        tmp_V_55_fu_790 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd54))) begin
        tmp_V_56_fu_794 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd55))) begin
        tmp_V_57_fu_798 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd56))) begin
        tmp_V_58_fu_802 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd57))) begin
        tmp_V_59_fu_806 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd3))) begin
        tmp_V_5_fu_590 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd58))) begin
        tmp_V_60_fu_810 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd59))) begin
        tmp_V_61_fu_814 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd60))) begin
        tmp_V_62_fu_818 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd61))) begin
        tmp_V_63_fu_822 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd62))) begin
        tmp_V_64_fu_826 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd63))) begin
        tmp_V_65_fu_830 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd64))) begin
        tmp_V_66_fu_834 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd65))) begin
        tmp_V_67_fu_838 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd66))) begin
        tmp_V_68_fu_842 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd67))) begin
        tmp_V_69_fu_846 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd4))) begin
        tmp_V_6_fu_594 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd68))) begin
        tmp_V_70_fu_850 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd69))) begin
        tmp_V_71_fu_854 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd70))) begin
        tmp_V_72_fu_858 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd71))) begin
        tmp_V_73_fu_862 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd72))) begin
        tmp_V_74_fu_866 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd73))) begin
        tmp_V_75_fu_870 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd74))) begin
        tmp_V_76_fu_874 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd75))) begin
        tmp_V_77_fu_878 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd76))) begin
        tmp_V_78_fu_882 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd77))) begin
        tmp_V_79_fu_886 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd5))) begin
        tmp_V_7_fu_598 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd78))) begin
        tmp_V_80_fu_890 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd79))) begin
        tmp_V_81_fu_894 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd80))) begin
        tmp_V_82_fu_898 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd81))) begin
        tmp_V_83_fu_902 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd82))) begin
        tmp_V_84_fu_906 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd83))) begin
        tmp_V_85_fu_910 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd84))) begin
        tmp_V_86_fu_914 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd85))) begin
        tmp_V_87_fu_918 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd86))) begin
        tmp_V_88_fu_922 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd87))) begin
        tmp_V_89_fu_926 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd6))) begin
        tmp_V_8_fu_602 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd88))) begin
        tmp_V_90_fu_930 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd89))) begin
        tmp_V_91_fu_934 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd90))) begin
        tmp_V_92_fu_938 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd91))) begin
        tmp_V_93_fu_942 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd92))) begin
        tmp_V_94_fu_946 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd93))) begin
        tmp_V_95_fu_950 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd94))) begin
        tmp_V_96_fu_954 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd95))) begin
        tmp_V_97_fu_958 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd96))) begin
        tmp_V_98_fu_962 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd97))) begin
        tmp_V_99_fu_966 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_3479_p1 == 8'd7))) begin
        tmp_V_9_fu_606 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_fu_570 <= tmp_V_260_fu_4871_p2;
    end
end

always @ (*) begin
    if ((icmp_ln248_fu_2165_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_6766 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_sig_allocacmp_nf_2_load = nf_3_fu_4898_p3;
    end else begin
        ap_sig_allocacmp_nf_2_load = nf_2_fu_1602;
    end
end

always @ (*) begin
    if (((icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op540_read_state2 == 1'b1))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_6766 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_6766 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln248_fu_2165_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TDATA_blk_n = weight_V_V_TVALID;
    end else begin
        weight_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_2165_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TREADY = 1'b1;
    end else begin
        weight_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((icmp_ln248_fu_2165_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((icmp_ln248_fu_2165_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln700_fu_4861_p2 = ($signed(sext_ln700_fu_4857_p1) + $signed(sext_ln170_fu_4830_p1));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op540_read_state2 == 1'b1)) | ((icmp_ln248_fu_2165_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op540_read_state2 == 1'b1)) | ((icmp_ln248_fu_2165_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op540_read_state2 == 1'b1)) | ((icmp_ln248_fu_2165_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op540_read_state2 == 1'b1)) | ((icmp_ln248_fu_2165_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)));
end

always @ (*) begin
    ap_block_state3_io = ((icmp_ln289_reg_6766 == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_reg_pp0_iter0_act_m_val_V_reg_1636 = 'bx;

always @ (*) begin
    ap_predicate_op540_read_state2 = ((icmp_ln252_fu_2180_p2 == 1'd1) & (icmp_ln248_fu_2165_p2 == 1'd0));
end

assign arg_V_read_assign_1_fu_4834_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1636[7:4]}};

assign i_fu_2171_p2 = (i_0_reg_1625 + 11'd1);

assign icmp_ln248_fu_2165_p2 = ((i_0_reg_1625 == 11'd1792) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_2180_p2 = ((ap_sig_allocacmp_nf_2_load == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln271_fu_4766_p2 = ((sf_1_fu_574 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln289_fu_4792_p2 = ((sf_fu_4786_p2 == 32'd256) ? 1'b1 : 1'b0);

assign icmp_ln301_fu_4892_p2 = ((nf_fu_4886_p2 == 32'd7) ? 1'b1 : 1'b0);

assign inElem_V_1_fu_2961_p257 = sf_1_fu_574[7:0];

assign nf_3_fu_4898_p3 = ((icmp_ln301_fu_4892_p2[0:0] === 1'b1) ? 32'd0 : nf_fu_4886_p2);

assign nf_fu_4886_p2 = (nf_2_fu_1602 + 32'd1);

assign out_V_V_TDATA = ($signed(res_V_fu_4806_p3) + $signed(sext_ln700_1_fu_4867_p1));

assign res_V_fu_4806_p3 = ((icmp_ln271_reg_6751[0:0] === 1'b1) ? 16'd0 : tmp_V_fu_570);

assign sext_ln170_fu_4830_p1 = mul_ln1352_fu_4824_p2;

assign sext_ln700_1_fu_4867_p1 = $signed(add_ln700_fu_4861_p2);

assign sext_ln700_fu_4857_p1 = mul_ln1352_1_fu_4851_p2;

assign sf_fu_4786_p2 = (32'd1 + sf_1_fu_574);

assign tmp_V_260_fu_4871_p2 = ($signed(res_V_fu_4806_p3) + $signed(sext_ln700_1_fu_4867_p1));

assign trunc_ln321_fu_3479_p1 = sf_1_fu_574[7:0];

assign trunc_ln647_1_fu_4813_p1 = ap_phi_reg_pp0_iter1_act_m_val_V_reg_1636[3:0];

assign trunc_ln647_fu_4772_p1 = weight_V_V_TDATA[3:0];

endmodule //StreamingFCLayer_Batch_6_Matrix_Vector_Activa
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActYie.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActYie_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActYie_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActYie(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActYie_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActYie_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbEo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcbEo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbEo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcbEo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcbEo_rom Thresholding_Batch_0_Thresholding_BatcbEo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/209a/hdl/memstream_singleblock.v

/*
 Copyright (c) 2020, Xilinx
 All rights reserved.

 Redistribution and use in source and binary forms, with or without
 modification, are permitted provided that the following conditions are met:

 * Redistributions of source code must retain the above copyright notice, this
   list of conditions and the following disclaimer.

 * Redistributions in binary form must reproduce the above copyright notice,
   this list of conditions and the following disclaimer in the documentation
   and/or other materials provided with the distribution.

 * Neither the name of FINN nor the names of its
   contributors may be used to endorse or promote products derived from
   this software without specific prior written permission.

 THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
 FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
 SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
 CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
 OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

/*
    Implements a lightweight streamer for up to 2 streams in a single block of memory
*/

module memstream_singleblock
#(
    parameter CONFIG_EN = 1,
    parameter NSTREAMS = 2,//1 up to 2

    parameter MEM_DEPTH = 512,
    parameter MEM_WIDTH = 32,
    parameter MEM_INIT = "./",
    parameter RAM_STYLE = "auto",

    //widths per stream
	parameter STRM0_WIDTH = 32,
	parameter STRM1_WIDTH = 32,

	//depths per stream
	parameter STRM0_DEPTH = 256,
	parameter STRM1_DEPTH = 256,

	//offsets for each stream
	parameter STRM0_OFFSET = 0,
	parameter STRM1_OFFSET = 256
)

(
    input aclk,
    input aresetn,

    //optional configuration interface compatible with ap_memory
	input [31:0] config_address,
	input config_ce,
	input config_we,
	input [MEM_WIDTH-1:0] config_d0,
	output [MEM_WIDTH-1:0] config_q0,
    output config_rack,

    //multiple output AXI Streams, TDATA width rounded to multiple of 8 bits
    input m_axis_0_tready,
    output m_axis_0_tvalid,
    output [((STRM0_WIDTH+7)/8)*8-1:0] m_axis_0_tdata,

    input m_axis_1_tready,
    output m_axis_1_tvalid,
    output [((STRM1_WIDTH+7)/8)*8-1:0] m_axis_1_tdata

);


//TODO: check that memory width is equal to the widest stream
//TODO: check that the stream depths and offsets make sense, and that the memory depth is sufficient (or calculate depth here?)
initial begin
    if((NSTREAMS < 1) | (NSTREAMS > 2)) begin
        $display("Invalid setting for NSTREAMS, please set in range [1,2]");
        $finish();
    end
end

//invert reset
wire rst;
assign rst = ~aresetn;

wire strm0_incr_en;
wire strm1_incr_en;

assign strm0_incr_en = m_axis_0_tready | ~m_axis_0_tvalid;
assign strm1_incr_en = m_axis_1_tready | ~m_axis_1_tvalid;

reg rack_shift[1:0];

generate
if(MEM_DEPTH > 1) begin: use_ram

//calculate width of memory address, with a minimum of 1 bit
localparam BLOCKADRWIDTH = $clog2(MEM_DEPTH);

reg [BLOCKADRWIDTH-1:0] strm0_addr = STRM0_OFFSET;
wire strm0_rst;
assign strm0_rst = strm0_incr_en & (strm0_addr == (STRM0_OFFSET + STRM0_DEPTH-1));

//one address counter per stream; more LUTs but keeps routing short and local
always @(posedge aclk) begin
    if(strm0_rst | rst)
        strm0_addr <= STRM0_OFFSET;
    else if(strm0_incr_en)
        strm0_addr <= strm0_addr + 1;
end

if(NSTREAMS == 1) begin: sdp

ramb18_sdp
#(
    .ID(0),
	.DWIDTH(MEM_WIDTH),
	.AWIDTH(BLOCKADRWIDTH),
    .DEPTH(MEM_DEPTH),
	.MEM_INIT(MEM_INIT),
    .RAM_STYLE(RAM_STYLE)
)
ram
(
	.clk(aclk),

    .ena(config_ce),
	.wea(config_we),
	.addra(config_address[BLOCKADRWIDTH-1:0]),
    .wdataa(config_d0),

    .enb(strm0_incr_en | config_ce),
    .enqb(strm0_incr_en | rack_shift[0]),
	.addrb(config_ce ? config_address[BLOCKADRWIDTH-1:0] : strm0_addr),
	.rdqb(m_axis_0_tdata)
);


end else begin: tdp

reg [BLOCKADRWIDTH-1:0] strm1_addr = STRM1_OFFSET;
wire strm1_rst;
assign strm1_rst = strm1_incr_en & (strm1_addr == (STRM1_OFFSET + STRM1_DEPTH-1));

always @(posedge aclk) begin
    if(strm1_rst | rst)
        strm1_addr <= STRM1_OFFSET;
    else if(strm1_incr_en)
        strm1_addr <= strm1_addr + 1;
end

ramb18_wf_dualport
#(
    .ID(0),
	.DWIDTH(MEM_WIDTH),
	.AWIDTH(BLOCKADRWIDTH),
    .DEPTH(MEM_DEPTH),
	.MEM_INIT(MEM_INIT),
    .RAM_STYLE(RAM_STYLE)
)
ram
(
	.clk(aclk),

	.wea(config_we),
    .ena(strm0_incr_en | config_ce),
    .enqa(strm0_incr_en | config_ce_r),
	.addra(config_we ? config_address[BLOCKADRWIDTH-1:0] : strm0_addr),
	.wdataa(config_d0),
	.rdqa(m_axis_0_tdata),

	.web(1'b0),
    .enb(strm1_incr_en),
    .enqb(strm1_incr_en),
	.addrb(strm1_addr),
	.wdatab('d0),
	.rdqb(m_axis_1_tdata)
);

end

end else begin: bypass

reg [MEM_WIDTH-1:0] singleval[0:0];
initial begin
    $readmemh({MEM_INIT,"memblock_0.dat"}, singleval, 0, 0);
end

always @(posedge aclk)
    if(config_ce & config_we)
        singleval[0] <= config_d0;

assign m_axis_0_tdata = singleval[0];
assign m_axis_1_tdata = singleval[0];

end
endgenerate

//signal valid after 2 tready cycles after initialization
//then stay valid
reg [1:0] tvalid_pipe0 = 2'd0;
reg [1:0] tvalid_pipe1 = 2'd0;

assign m_axis_0_tvalid = tvalid_pipe0[1];
assign m_axis_1_tvalid = tvalid_pipe1[1];

always @(posedge aclk) begin
    if(rst) begin
        tvalid_pipe0 <= 0;
    end else if(strm0_incr_en) begin
        tvalid_pipe0[0] <= 1;
        tvalid_pipe0[1] <= tvalid_pipe0[0];
    end
end

always @(posedge aclk) begin
    if(rst) begin
        tvalid_pipe1 <= 0;
    end else if(strm1_incr_en) begin
        tvalid_pipe1[0] <= 1;
        tvalid_pipe1[1] <= tvalid_pipe1[0];
    end
end

always @(posedge aclk) begin
    rack_shift[0] <= config_ce & ~config_we;
    rack_shift[1] <= rack_shift[0];
end

assign config_rack = rack_shift[1];
assign config_q0 = m_axis_0_tdata;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Act0iy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Act0iy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Act0iy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Act0iy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Act0iy_rom StreamingFCLayer_Batch_1_Matrix_Vector_Act0iy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActNgs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActNgs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActNgs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActNgs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActNgs_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActNgs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActFfa.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActFfa_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActFfa_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActFfa(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActFfa_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActFfa_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/regslice_core.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module regslice_both
#(parameter 
    DataWidth=32
)(
    input ap_clk ,
    input ap_rst,

    input [DataWidth-1:0] data_in , 
    input vld_in , 
    output ack_in ,
    output [DataWidth-1:0] data_out, 
    output vld_out,
    input ack_out,
    output apdone_blk
);
 
localparam W = DataWidth+1;

wire [W-1:0] cdata;
wire cstop;
wire [W-1:0] idata;
wire istop;
wire [W-1:0] odata;
wire ostop;

reg [1:0] count;

ibuf #(
  .W(W)
)
ibuf_inst(
  .clk(ap_clk),
  .reset(ap_rst),
  .idata(idata),
  .istop(istop),
  .cdata(cdata),
  .cstop(cstop)
);
 
 
obuf #(
  .W(W)
)
obuf_inst(
  .clk(ap_clk),
  .reset(ap_rst),
  .cdata(cdata),
  .cstop(cstop),
  .odata(odata),
  .ostop(ostop)
);

assign idata = {vld_in, data_in};
assign ack_in = ~istop;

assign vld_out = odata[W-1];
assign data_out = odata[W-2:0];
assign ostop = ~ack_out;

// count, indicate how many data in the regslice.
// 00 - null
// 10 - 0
// 11 - 1
// 01 - 2
always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        count <= 2'd0;
    end else begin
        if ((((2'd2 == count) & (1'b0 == vld_in)) | ((2'd3 == count) & (1'b0 == vld_in) & (1'b1 == ack_out)))) begin
            count <= 2'd2;
        end else if ((((2'd1 == count) & (1'b0 == ack_out)) | ((2'd3 == count) & (1'b0 == ack_out) & (1'b1 == vld_in)))) begin
            count <= 2'd1;
        end else if (((~((1'b0 == vld_in) & (1'b1 == ack_out)) & ~((1'b0 == ack_out) & (1'b1 == vld_in)) & (2'd3 == count)) | ((2'd1 == count) & (1'b1 == ack_out)) | ((2'd2 == count) & (1'b1 == vld_in)))) begin
            count <= 2'd3;
        end else begin
            count <= 2'd2;
        end
    end
end

assign apdone_blk = ((count == 2'd3 && ack_out == 1'b0) | (count == 2'd1));

endmodule // both


module regslice_forward 
#(parameter 
    DataWidth=32
)(
    input ap_clk ,
    input ap_rst,

    input [DataWidth-1:0] data_in , 
    input vld_in , 
    output ack_in ,
    output [DataWidth-1:0] data_out, 
    output vld_out,
    input ack_out,
    output apdone_blk
);
 
localparam W = DataWidth+1;

wire [W-1:0] cdata;
wire cstop;
wire [W-1:0] idata;
wire istop;
wire [W-1:0] odata;
wire ostop;

obuf #(
  .W(W)
)
obuf_inst(
  .clk(ap_clk),
  .reset(ap_rst),
  .cdata(idata),
  .cstop(istop),
  .odata(odata),
  .ostop(ostop)
);

assign idata = {vld_in, data_in};
assign ack_in = ~istop;

assign vld_out = odata[W-1];
assign data_out = odata[W-2:0];
assign ostop = ~ack_out;

assign apdone_blk = ((ap_rst == 1'b0)&(1'b0 == ack_out)&(1'b1 == vld_out));

endmodule //forward


module regslice_reverse 
#(parameter 
    DataWidth=32
)(
    input ap_clk ,
    input ap_rst,

    input [DataWidth-1:0] data_in , 
    input vld_in , 
    output ack_in ,
    output [DataWidth-1:0] data_out, 
    output vld_out,
    input ack_out,
    output apdone_blk
);
 
localparam W = DataWidth+1;

wire [W-1:0] cdata;
wire cstop;
wire [W-1:0] idata;
wire istop;
wire [W-1:0] odata;
wire ostop;

ibuf #(
  .W(W)
)
ibuf_inst(
  .clk(ap_clk),
  .reset(ap_rst),
  .idata(idata),
  .istop(istop),
  .cdata(odata),
  .cstop(ostop)
);
 
assign idata = {vld_in, data_in};
assign ack_in = ~istop;

assign vld_out = odata[W-1];
assign data_out = odata[W-2:0];
assign ostop = ~ack_out;

assign apdone_blk = ((ap_rst == 1'b0)&(ack_in == 1'b0));

endmodule //reverse

module regslice_both_w1 
#(parameter 
    DataWidth=32
)(
    input ap_clk ,
    input ap_rst,

    input data_in , 
    input vld_in , 
    output ack_in ,
    output data_out, 
    output vld_out,
    input ack_out,
    output apdone_blk
);
 
localparam W = 2;

wire [W-1:0] cdata;
wire cstop;
wire [W-1:0] idata;
wire istop;
wire [W-1:0] odata;
wire ostop;

reg [1:0] count;

ibuf #(
  .W(W)
)
ibuf_inst(
  .clk(ap_clk),
  .reset(ap_rst),
  .idata(idata),
  .istop(istop),
  .cdata(cdata),
  .cstop(cstop)
);
 
 
obuf #(
  .W(W)
)
obuf_inst(
  .clk(ap_clk),
  .reset(ap_rst),
  .cdata(cdata),
  .cstop(cstop),
  .odata(odata),
  .ostop(ostop)
);

assign idata = {vld_in, data_in};
assign ack_in = ~istop;

assign vld_out = odata[W-1];
assign data_out = odata[W-2:0];
assign ostop = ~ack_out;
// count, indicate how many data in the regslice.
// 00 - null
// 10 - 0
// 11 - 1
// 01 - 2
always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        count <= 2'd0;
    end else begin
        if ((((2'd2 == count) & (1'b0 == vld_in)) | ((2'd3 == count) & (1'b0 == vld_in) & (1'b1 == ack_out)))) begin
            count <= 2'd2;
        end else if ((((2'd1 == count) & (1'b0 == ack_out)) | ((2'd3 == count) & (1'b0 == ack_out) & (1'b1 == vld_in)))) begin
            count <= 2'd1;
        end else if (((~((1'b0 == vld_in) & (1'b1 == ack_out)) & ~((1'b0 == ack_out) & (1'b1 == vld_in)) & (2'd3 == count)) | ((2'd1 == count) & (1'b1 == ack_out)) | ((2'd2 == count) & (1'b1 == vld_in)))) begin
            count <= 2'd3;
        end else begin
            count <= 2'd2;
        end
    end
end

assign apdone_blk = ((count == 2'd3 && ack_out == 1'b0) | (count == 2'd1));

endmodule // both


module regslice_forward_w1 
#(parameter 
    DataWidth=1
)(
    input ap_clk ,
    input ap_rst,

    input data_in , 
    input vld_in , 
    output ack_in ,
    output data_out, 
    output vld_out,
    input ack_out,
    output apdone_blk
);
 
localparam W = 2;

wire [W-1:0] cdata;
wire cstop;
wire [W-1:0] idata;
wire istop;
wire [W-1:0] odata;
wire ostop;

obuf #(
  .W(W)
)
obuf_inst(
  .clk(ap_clk),
  .reset(ap_rst),
  .cdata(idata),
  .cstop(istop),
  .odata(odata),
  .ostop(ostop)
);

assign idata = {vld_in, data_in};
assign ack_in = ~istop;

assign vld_out = odata[W-1];
assign data_out = odata[W-2:0];
assign ostop = ~ack_out;

assign apdone_blk = ((ap_rst == 1'b0)&(1'b0 == ack_out)&(1'b1 == vld_out));

endmodule //forward


module regslice_reverse_w1 
#(parameter 
    DataWidth=1
)(
    input ap_clk ,
    input ap_rst,

    input data_in , 
    input vld_in , 
    output ack_in ,
    output data_out, 
    output vld_out,
    input ack_out,
    output apdone_blk
);
 
localparam W = 2;

wire [W-1:0] cdata;
wire cstop;
wire [W-1:0] idata;
wire istop;
wire [W-1:0] odata;
wire ostop;

ibuf #(
  .W(W)
)
ibuf_inst(
  .clk(ap_clk),
  .reset(ap_rst),
  .idata(idata),
  .istop(istop),
  .cdata(odata),
  .cstop(ostop)
);
 
assign idata = {vld_in, data_in};
assign ack_in = ~istop;

assign vld_out = odata[W-1];
assign data_out = odata[W-2:0];
assign ostop = ~ack_out;

assign apdone_blk = ((ap_rst == 1'b0)&(ack_in == 1'b0));

endmodule //reverse


module ibuf 
#(
    parameter W=32
)(
    input clk ,
    input reset,
    input [W-1:0] idata, 
    output istop ,
    output [W-1:0] cdata, 
    input cstop 
);
 
reg [W-1:0] ireg = {1'b0, {{W-1}{1'b0}}}; // Empty
 
assign istop = reset ? 1'b1 : ireg[W-1]; // Stop if buffering
assign cdata = istop ? ireg : idata ; // Send buffered
 
always @(posedge clk)
    if(reset)
        ireg <= {1'b0, {{W-1}{1'b0}}}; // Empty 
    else begin
        if (!cstop && ireg [W-1]) // Will core consume?
            ireg <= {1'b0, {{W-1}{1'b0}}}; // Yes: empty buffer
        else if ( cstop && !ireg[W-1]) // Core stop, empty?
            ireg <= idata; // Yes: load buffer
    end
 
endmodule

// Forward mode
module obuf 
#(
    parameter W=32
)(
    input clk ,
    input reset,
    input [W-1:0] cdata ,
    output cstop ,
    output reg [W-1:0] odata,
    input ostop 
);

// Stop the core when buffer full and output not ready
assign cstop = reset? 1'b1 : (odata[W-1] & ostop);
 
always @(posedge clk)
    if(reset)
        odata <= {1'b0, {{W-1}{1'b0}}};
    else
        if (!cstop) begin// Can we accept more data?
            odata <= cdata; // Yes: load the buffer
        end

endmodule

    
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Act2iS.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Act2iS_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Act2iS_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Act2iS(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Act2iS_rom StreamingFCLayer_Batch_1_Matrix_Vector_Act2iS_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActMgi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActMgi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActMgi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActMgi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActMgi_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActMgi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actncg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actncg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actncg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actncg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actncg_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actncg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbsm.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbsm_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbsm_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbsm(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbsm_rom Thresholding_Batch_0_Thresholding_Batcbsm_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActxdS.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActxdS_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActxdS_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActxdS(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActxdS_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActxdS_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_BatclbW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_BatclbW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_BatclbW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_BatclbW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_BatclbW_rom Thresholding_Batch_1_Thresholding_BatclbW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/c3f7/hdl/verilog/LabelSelect_Batch_0_LabelSelect_Batch.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module LabelSelect_Batch_0_LabelSelect_Batch (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_state2 = 3'd2;
parameter    ap_ST_fsm_state3 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [15:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln374_fu_83_p2;
reg    out_V_V_TDATA_blk_n;
wire    ap_CS_fsm_state3;
wire   [2:0] add_ln397_fu_89_p2;
reg    ap_block_state2;
wire   [15:0] topval_0_V_1_fu_105_p3;
reg   [15:0] topval_V_0_0_reg_57;
reg   [2:0] idx_0_0_reg_68;
reg   [7:0] tmp_V_fu_40;
wire   [7:0] toplabels_0_V_1_fu_113_p3;
wire   [0:0] icmp_ln895_fu_95_p2;
wire   [7:0] toplabels_0_V_fu_101_p1;
reg   [2:0] ap_NS_fsm;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if ((~((icmp_ln374_fu_83_p2 == 1'd0) & (in_V_V_TVALID == 1'b0)) & (icmp_ln374_fu_83_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        idx_0_0_reg_68 <= add_ln397_fu_89_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        idx_0_0_reg_68 <= 3'd0;
    end
end

always @ (posedge ap_clk) begin
    if ((~((icmp_ln374_fu_83_p2 == 1'd0) & (in_V_V_TVALID == 1'b0)) & (icmp_ln374_fu_83_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        topval_V_0_0_reg_57 <= topval_0_V_1_fu_105_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        topval_V_0_0_reg_57 <= 16'd32768;
    end
end

always @ (posedge ap_clk) begin
    if ((~((icmp_ln374_fu_83_p2 == 1'd0) & (in_V_V_TVALID == 1'b0)) & (icmp_ln374_fu_83_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        tmp_V_fu_40 <= toplabels_0_V_1_fu_113_p3;
    end
end

always @ (*) begin
    if ((((out_V_V_TREADY == 1'b1) & (1'b1 == ap_CS_fsm_state3)) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((out_V_V_TREADY == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln374_fu_83_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((icmp_ln374_fu_83_p2 == 1'd0) & (in_V_V_TVALID == 1'b0)) & (icmp_ln374_fu_83_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((out_V_V_TREADY == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if ((~((icmp_ln374_fu_83_p2 == 1'd0) & (in_V_V_TVALID == 1'b0)) & (icmp_ln374_fu_83_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else if ((~((icmp_ln374_fu_83_p2 == 1'd0) & (in_V_V_TVALID == 1'b0)) & (icmp_ln374_fu_83_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end
        end
        ap_ST_fsm_state3 : begin
            if (((out_V_V_TREADY == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln397_fu_89_p2 = (idx_0_0_reg_68 + 3'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

always @ (*) begin
    ap_block_state2 = ((icmp_ln374_fu_83_p2 == 1'd0) & (in_V_V_TVALID == 1'b0));
end

assign icmp_ln374_fu_83_p2 = ((idx_0_0_reg_68 == 3'd7) ? 1'b1 : 1'b0);

assign icmp_ln895_fu_95_p2 = (($signed(in_V_V_TDATA) > $signed(topval_V_0_0_reg_57)) ? 1'b1 : 1'b0);

assign out_V_V_TDATA = tmp_V_fu_40;

assign toplabels_0_V_1_fu_113_p3 = ((icmp_ln895_fu_95_p2[0:0] === 1'b1) ? toplabels_0_V_fu_101_p1 : tmp_V_fu_40);

assign toplabels_0_V_fu_101_p1 = idx_0_0_reg_68;

assign topval_0_V_1_fu_105_p3 = ((icmp_ln895_fu_95_p2[0:0] === 1'b1) ? in_V_V_TDATA : topval_V_0_0_reg_57);

endmodule //LabelSelect_Batch_0_LabelSelect_Batch
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbGp.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcbGp_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbGp_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcbGp(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcbGp_rom Thresholding_Batch_0_Thresholding_BatcbGp_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActCeG.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActCeG_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActCeG_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActCeG(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActCeG_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActCeG_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActWhU.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActWhU_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActWhU_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActWhU(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActWhU_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActWhU_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActjbC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActjbC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActjbC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActjbC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActjbC_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActjbC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_6_0/synth/finn_design_StreamingFCLayer_Batch_6_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFCLayer_Batch_6:1.0
// IP Revision: 2101301316

(* X_CORE_INFO = "StreamingFCLayer_Batch_6_StreamingFCLayer_Batch_6,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_6_0,StreamingFCLayer_Batch_6_StreamingFCLayer_Batch_6,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_6_0,StreamingFCLayer_Batch_6_StreamingFCLayer_Batch_6,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFCLayer_Batch_6,x_ipVersion=1.0,x_ipCoreRevision=2101301316,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_6_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  weights_V_V_TVALID,
  weights_V_V_TREADY,
  weights_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:weights_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [7 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TVALID" *)
input wire weights_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TREADY" *)
output wire weights_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME weights_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TDATA" *)
input wire [7 : 0] weights_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;

  StreamingFCLayer_Batch_6_StreamingFCLayer_Batch_6 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .weights_V_V_TVALID(weights_V_V_TVALID),
    .weights_V_V_TREADY(weights_V_V_TREADY),
    .weights_V_V_TDATA(weights_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_ConvolutionInputGenerator_0_0/synth/finn_design_ConvolutionInputGenerator_0_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:ConvolutionInputGenerator_0:1.0
// IP Revision: 2101301318

(* X_CORE_INFO = "ConvolutionInputGenerator_0_ConvolutionInputGenerator_0,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_ConvolutionInputGenerator_0_0,ConvolutionInputGenerator_0_ConvolutionInputGenerator_0,{}" *)
(* CORE_GENERATION_INFO = "finn_design_ConvolutionInputGenerator_0_0,ConvolutionInputGenerator_0_ConvolutionInputGenerator_0,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=ConvolutionInputGenerator_0,x_ipVersion=1.0,x_ipCoreRevision=2101301318,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_ConvolutionInputGenerator_0_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [7 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;

  ConvolutionInputGenerator_0_ConvolutionInputGenerator_0 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actncg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actncg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actncg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actncg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actncg_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actncg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_12_0/synth/finn_design_StreamingFIFO_12_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_12:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_12,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_12_0,StreamingFIFO_12,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_12_0,StreamingFIFO_12,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_12,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_12_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [31 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 4, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [31 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 4, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_12 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActjbC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActjbC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActjbC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActjbC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActjbC_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActjbC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_Thresholding_Batch_0_0/synth/finn_design_Thresholding_Batch_0_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:Thresholding_Batch_0:1.0
// IP Revision: 2101301319

(* X_CORE_INFO = "Thresholding_Batch_0_Thresholding_Batch_0,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_Thresholding_Batch_0_0,Thresholding_Batch_0_Thresholding_Batch_0,{}" *)
(* CORE_GENERATION_INFO = "finn_design_Thresholding_Batch_0_0,Thresholding_Batch_0_Thresholding_Batch_0,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=Thresholding_Batch_0,x_ipVersion=1.0,x_ipCoreRevision=2101301319,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_Thresholding_Batch_0_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [7 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;

  Thresholding_Batch_0_Thresholding_Batch_0 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_Thresholding_Batch_2_0/synth/finn_design_Thresholding_Batch_2_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:Thresholding_Batch_2:1.0
// IP Revision: 2101301315

(* X_CORE_INFO = "Thresholding_Batch_2_Thresholding_Batch_2,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_Thresholding_Batch_2_0,Thresholding_Batch_2_Thresholding_Batch_2,{}" *)
(* CORE_GENERATION_INFO = "finn_design_Thresholding_Batch_2_0,Thresholding_Batch_2_Thresholding_Batch_2,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=Thresholding_Batch_2,x_ipVersion=1.0,x_ipCoreRevision=2101301315,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_Thresholding_Batch_2_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;

  Thresholding_Batch_2_Thresholding_Batch_2 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActRg6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActRg6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActRg6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActRg6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActRg6_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActRg6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatclbW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatclbW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 4;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatclbW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatclbW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd4;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatclbW_rom Thresholding_Batch_0_Thresholding_BatclbW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccCy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccCy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccCy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccCy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccCy_rom Thresholding_Batch_0_Thresholding_BatccCy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batch.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module Thresholding_Batch_0_Thresholding_Batch (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state6 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [7:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [1:0] threshs_m_thresholds_254_address0;
reg    threshs_m_thresholds_254_ce0;
wire   [0:0] threshs_m_thresholds_254_q0;
wire   [1:0] threshs_m_thresholds_253_address0;
reg    threshs_m_thresholds_253_ce0;
wire   [1:0] threshs_m_thresholds_253_q0;
wire   [1:0] threshs_m_thresholds_142_address0;
reg    threshs_m_thresholds_142_ce0;
wire   [0:0] threshs_m_thresholds_142_q0;
wire   [1:0] threshs_m_thresholds_76_address0;
reg    threshs_m_thresholds_76_ce0;
wire   [2:0] threshs_m_thresholds_76_q0;
wire   [1:0] threshs_m_thresholds_65_address0;
reg    threshs_m_thresholds_65_ce0;
wire   [2:0] threshs_m_thresholds_65_q0;
wire   [1:0] threshs_m_thresholds_54_address0;
reg    threshs_m_thresholds_54_ce0;
wire   [1:0] threshs_m_thresholds_54_q0;
wire   [1:0] threshs_m_thresholds_43_address0;
reg    threshs_m_thresholds_43_ce0;
wire   [0:0] threshs_m_thresholds_43_q0;
wire   [1:0] threshs_m_thresholds_32_address0;
reg    threshs_m_thresholds_32_ce0;
wire   [3:0] threshs_m_thresholds_32_q0;
wire   [1:0] threshs_m_thresholds_21_address0;
reg    threshs_m_thresholds_21_ce0;
wire   [3:0] threshs_m_thresholds_21_q0;
wire   [1:0] threshs_m_thresholds_10_address0;
reg    threshs_m_thresholds_10_ce0;
wire   [3:0] threshs_m_thresholds_10_q0;
wire   [1:0] threshs_m_thresholds_252_address0;
reg    threshs_m_thresholds_252_ce0;
wire   [3:0] threshs_m_thresholds_252_q0;
wire   [1:0] threshs_m_thresholds_241_address0;
reg    threshs_m_thresholds_241_ce0;
wire   [2:0] threshs_m_thresholds_241_q0;
wire   [1:0] threshs_m_thresholds_230_address0;
reg    threshs_m_thresholds_230_ce0;
wire   [2:0] threshs_m_thresholds_230_q0;
wire   [1:0] threshs_m_thresholds_219_address0;
reg    threshs_m_thresholds_219_ce0;
wire   [1:0] threshs_m_thresholds_219_q0;
wire   [1:0] threshs_m_thresholds_208_address0;
reg    threshs_m_thresholds_208_ce0;
wire   [0:0] threshs_m_thresholds_208_q0;
wire   [1:0] threshs_m_thresholds_197_address0;
reg    threshs_m_thresholds_197_ce0;
wire   [4:0] threshs_m_thresholds_197_q0;
wire   [1:0] threshs_m_thresholds_186_address0;
reg    threshs_m_thresholds_186_ce0;
wire   [4:0] threshs_m_thresholds_186_q0;
wire   [1:0] threshs_m_thresholds_175_address0;
reg    threshs_m_thresholds_175_ce0;
wire   [4:0] threshs_m_thresholds_175_q0;
wire   [1:0] threshs_m_thresholds_164_address0;
reg    threshs_m_thresholds_164_ce0;
wire   [4:0] threshs_m_thresholds_164_q0;
wire   [1:0] threshs_m_thresholds_153_address0;
reg    threshs_m_thresholds_153_ce0;
wire   [4:0] threshs_m_thresholds_153_q0;
wire   [1:0] threshs_m_thresholds_141_address0;
reg    threshs_m_thresholds_141_ce0;
wire   [4:0] threshs_m_thresholds_141_q0;
wire   [1:0] threshs_m_thresholds_130_address0;
reg    threshs_m_thresholds_130_ce0;
wire   [4:0] threshs_m_thresholds_130_q0;
wire   [1:0] threshs_m_thresholds_119_address0;
reg    threshs_m_thresholds_119_ce0;
wire   [4:0] threshs_m_thresholds_119_q0;
wire   [1:0] threshs_m_thresholds_108_address0;
reg    threshs_m_thresholds_108_ce0;
wire   [3:0] threshs_m_thresholds_108_q0;
wire   [1:0] threshs_m_thresholds_97_address0;
reg    threshs_m_thresholds_97_ce0;
wire   [3:0] threshs_m_thresholds_97_q0;
wire   [1:0] threshs_m_thresholds_86_address0;
reg    threshs_m_thresholds_86_ce0;
wire   [3:0] threshs_m_thresholds_86_q0;
wire   [1:0] threshs_m_thresholds_80_address0;
reg    threshs_m_thresholds_80_ce0;
wire   [3:0] threshs_m_thresholds_80_q0;
wire   [1:0] threshs_m_thresholds_79_address0;
reg    threshs_m_thresholds_79_ce0;
wire   [2:0] threshs_m_thresholds_79_q0;
wire   [1:0] threshs_m_thresholds_78_address0;
reg    threshs_m_thresholds_78_ce0;
wire   [2:0] threshs_m_thresholds_78_q0;
wire   [1:0] threshs_m_thresholds_77_address0;
reg    threshs_m_thresholds_77_ce0;
wire   [1:0] threshs_m_thresholds_77_q0;
wire   [1:0] threshs_m_thresholds_75_address0;
reg    threshs_m_thresholds_75_ce0;
wire   [0:0] threshs_m_thresholds_75_q0;
wire   [1:0] threshs_m_thresholds_74_address0;
reg    threshs_m_thresholds_74_ce0;
wire   [5:0] threshs_m_thresholds_74_q0;
wire   [1:0] threshs_m_thresholds_73_address0;
reg    threshs_m_thresholds_73_ce0;
wire   [5:0] threshs_m_thresholds_73_q0;
wire   [1:0] threshs_m_thresholds_72_address0;
reg    threshs_m_thresholds_72_ce0;
wire   [5:0] threshs_m_thresholds_72_q0;
wire   [1:0] threshs_m_thresholds_71_address0;
reg    threshs_m_thresholds_71_ce0;
wire   [5:0] threshs_m_thresholds_71_q0;
wire   [1:0] threshs_m_thresholds_70_address0;
reg    threshs_m_thresholds_70_ce0;
wire   [5:0] threshs_m_thresholds_70_q0;
wire   [1:0] threshs_m_thresholds_69_address0;
reg    threshs_m_thresholds_69_ce0;
wire   [5:0] threshs_m_thresholds_69_q0;
wire   [1:0] threshs_m_thresholds_68_address0;
reg    threshs_m_thresholds_68_ce0;
wire   [5:0] threshs_m_thresholds_68_q0;
wire   [1:0] threshs_m_thresholds_67_address0;
reg    threshs_m_thresholds_67_ce0;
wire   [5:0] threshs_m_thresholds_67_q0;
wire   [1:0] threshs_m_thresholds_66_address0;
reg    threshs_m_thresholds_66_ce0;
wire   [5:0] threshs_m_thresholds_66_q0;
wire   [1:0] threshs_m_thresholds_64_address0;
reg    threshs_m_thresholds_64_ce0;
wire   [5:0] threshs_m_thresholds_64_q0;
wire   [1:0] threshs_m_thresholds_63_address0;
reg    threshs_m_thresholds_63_ce0;
wire   [5:0] threshs_m_thresholds_63_q0;
wire   [1:0] threshs_m_thresholds_62_address0;
reg    threshs_m_thresholds_62_ce0;
wire   [5:0] threshs_m_thresholds_62_q0;
wire   [1:0] threshs_m_thresholds_61_address0;
reg    threshs_m_thresholds_61_ce0;
wire   [5:0] threshs_m_thresholds_61_q0;
wire   [1:0] threshs_m_thresholds_60_address0;
reg    threshs_m_thresholds_60_ce0;
wire   [5:0] threshs_m_thresholds_60_q0;
wire   [1:0] threshs_m_thresholds_59_address0;
reg    threshs_m_thresholds_59_ce0;
wire   [5:0] threshs_m_thresholds_59_q0;
wire   [1:0] threshs_m_thresholds_58_address0;
reg    threshs_m_thresholds_58_ce0;
wire   [5:0] threshs_m_thresholds_58_q0;
wire   [1:0] threshs_m_thresholds_57_address0;
reg    threshs_m_thresholds_57_ce0;
wire   [4:0] threshs_m_thresholds_57_q0;
wire   [1:0] threshs_m_thresholds_56_address0;
reg    threshs_m_thresholds_56_ce0;
wire   [4:0] threshs_m_thresholds_56_q0;
wire   [1:0] threshs_m_thresholds_55_address0;
reg    threshs_m_thresholds_55_ce0;
wire   [4:0] threshs_m_thresholds_55_q0;
wire   [1:0] threshs_m_thresholds_53_address0;
reg    threshs_m_thresholds_53_ce0;
wire   [4:0] threshs_m_thresholds_53_q0;
wire   [1:0] threshs_m_thresholds_52_address0;
reg    threshs_m_thresholds_52_ce0;
wire   [4:0] threshs_m_thresholds_52_q0;
wire   [1:0] threshs_m_thresholds_51_address0;
reg    threshs_m_thresholds_51_ce0;
wire   [4:0] threshs_m_thresholds_51_q0;
wire   [1:0] threshs_m_thresholds_50_address0;
reg    threshs_m_thresholds_50_ce0;
wire   [4:0] threshs_m_thresholds_50_q0;
wire   [1:0] threshs_m_thresholds_49_address0;
reg    threshs_m_thresholds_49_ce0;
wire   [4:0] threshs_m_thresholds_49_q0;
wire   [1:0] threshs_m_thresholds_48_address0;
reg    threshs_m_thresholds_48_ce0;
wire   [3:0] threshs_m_thresholds_48_q0;
wire   [1:0] threshs_m_thresholds_47_address0;
reg    threshs_m_thresholds_47_ce0;
wire   [3:0] threshs_m_thresholds_47_q0;
wire   [1:0] threshs_m_thresholds_46_address0;
reg    threshs_m_thresholds_46_ce0;
wire   [3:0] threshs_m_thresholds_46_q0;
wire   [1:0] threshs_m_thresholds_45_address0;
reg    threshs_m_thresholds_45_ce0;
wire   [3:0] threshs_m_thresholds_45_q0;
wire   [1:0] threshs_m_thresholds_44_address0;
reg    threshs_m_thresholds_44_ce0;
wire   [2:0] threshs_m_thresholds_44_q0;
wire   [1:0] threshs_m_thresholds_42_address0;
reg    threshs_m_thresholds_42_ce0;
wire   [2:0] threshs_m_thresholds_42_q0;
wire   [1:0] threshs_m_thresholds_41_address0;
reg    threshs_m_thresholds_41_ce0;
wire   [1:0] threshs_m_thresholds_41_q0;
wire   [1:0] threshs_m_thresholds_40_address0;
reg    threshs_m_thresholds_40_ce0;
wire   [0:0] threshs_m_thresholds_40_q0;
wire   [1:0] threshs_m_thresholds_39_address0;
reg    threshs_m_thresholds_39_ce0;
wire   [6:0] threshs_m_thresholds_39_q0;
wire   [1:0] threshs_m_thresholds_38_address0;
reg    threshs_m_thresholds_38_ce0;
wire   [6:0] threshs_m_thresholds_38_q0;
wire   [1:0] threshs_m_thresholds_37_address0;
reg    threshs_m_thresholds_37_ce0;
wire   [6:0] threshs_m_thresholds_37_q0;
wire   [1:0] threshs_m_thresholds_36_address0;
reg    threshs_m_thresholds_36_ce0;
wire   [6:0] threshs_m_thresholds_36_q0;
wire   [1:0] threshs_m_thresholds_35_address0;
reg    threshs_m_thresholds_35_ce0;
wire   [6:0] threshs_m_thresholds_35_q0;
wire   [1:0] threshs_m_thresholds_34_address0;
reg    threshs_m_thresholds_34_ce0;
wire   [6:0] threshs_m_thresholds_34_q0;
wire   [1:0] threshs_m_thresholds_33_address0;
reg    threshs_m_thresholds_33_ce0;
wire   [6:0] threshs_m_thresholds_33_q0;
wire   [1:0] threshs_m_thresholds_31_address0;
reg    threshs_m_thresholds_31_ce0;
wire   [6:0] threshs_m_thresholds_31_q0;
wire   [1:0] threshs_m_thresholds_30_address0;
reg    threshs_m_thresholds_30_ce0;
wire   [6:0] threshs_m_thresholds_30_q0;
wire   [1:0] threshs_m_thresholds_29_address0;
reg    threshs_m_thresholds_29_ce0;
wire   [6:0] threshs_m_thresholds_29_q0;
wire   [1:0] threshs_m_thresholds_28_address0;
reg    threshs_m_thresholds_28_ce0;
wire   [6:0] threshs_m_thresholds_28_q0;
wire   [1:0] threshs_m_thresholds_27_address0;
reg    threshs_m_thresholds_27_ce0;
wire   [6:0] threshs_m_thresholds_27_q0;
wire   [1:0] threshs_m_thresholds_26_address0;
reg    threshs_m_thresholds_26_ce0;
wire   [6:0] threshs_m_thresholds_26_q0;
wire   [1:0] threshs_m_thresholds_25_address0;
reg    threshs_m_thresholds_25_ce0;
wire   [6:0] threshs_m_thresholds_25_q0;
wire   [1:0] threshs_m_thresholds_24_address0;
reg    threshs_m_thresholds_24_ce0;
wire   [6:0] threshs_m_thresholds_24_q0;
wire   [1:0] threshs_m_thresholds_23_address0;
reg    threshs_m_thresholds_23_ce0;
wire   [6:0] threshs_m_thresholds_23_q0;
wire   [1:0] threshs_m_thresholds_22_address0;
reg    threshs_m_thresholds_22_ce0;
wire   [6:0] threshs_m_thresholds_22_q0;
wire   [1:0] threshs_m_thresholds_20_address0;
reg    threshs_m_thresholds_20_ce0;
wire   [6:0] threshs_m_thresholds_20_q0;
wire   [1:0] threshs_m_thresholds_19_address0;
reg    threshs_m_thresholds_19_ce0;
wire   [6:0] threshs_m_thresholds_19_q0;
wire   [1:0] threshs_m_thresholds_18_address0;
reg    threshs_m_thresholds_18_ce0;
wire   [6:0] threshs_m_thresholds_18_q0;
wire   [1:0] threshs_m_thresholds_17_address0;
reg    threshs_m_thresholds_17_ce0;
wire   [6:0] threshs_m_thresholds_17_q0;
wire   [1:0] threshs_m_thresholds_16_address0;
reg    threshs_m_thresholds_16_ce0;
wire   [6:0] threshs_m_thresholds_16_q0;
wire   [1:0] threshs_m_thresholds_15_address0;
reg    threshs_m_thresholds_15_ce0;
wire   [6:0] threshs_m_thresholds_15_q0;
wire   [1:0] threshs_m_thresholds_14_address0;
reg    threshs_m_thresholds_14_ce0;
wire   [6:0] threshs_m_thresholds_14_q0;
wire   [1:0] threshs_m_thresholds_13_address0;
reg    threshs_m_thresholds_13_ce0;
wire   [6:0] threshs_m_thresholds_13_q0;
wire   [1:0] threshs_m_thresholds_12_address0;
reg    threshs_m_thresholds_12_ce0;
wire   [6:0] threshs_m_thresholds_12_q0;
wire   [1:0] threshs_m_thresholds_11_address0;
reg    threshs_m_thresholds_11_ce0;
wire   [6:0] threshs_m_thresholds_11_q0;
wire   [1:0] threshs_m_thresholds_9_address0;
reg    threshs_m_thresholds_9_ce0;
wire   [6:0] threshs_m_thresholds_9_q0;
wire   [1:0] threshs_m_thresholds_8_address0;
reg    threshs_m_thresholds_8_ce0;
wire   [6:0] threshs_m_thresholds_8_q0;
wire   [1:0] threshs_m_thresholds_7_address0;
reg    threshs_m_thresholds_7_ce0;
wire   [6:0] threshs_m_thresholds_7_q0;
wire   [1:0] threshs_m_thresholds_6_address0;
reg    threshs_m_thresholds_6_ce0;
wire   [6:0] threshs_m_thresholds_6_q0;
wire   [1:0] threshs_m_thresholds_5_address0;
reg    threshs_m_thresholds_5_ce0;
wire   [6:0] threshs_m_thresholds_5_q0;
wire   [1:0] threshs_m_thresholds_4_address0;
reg    threshs_m_thresholds_4_ce0;
wire   [5:0] threshs_m_thresholds_4_q0;
wire   [1:0] threshs_m_thresholds_3_address0;
reg    threshs_m_thresholds_3_ce0;
wire   [5:0] threshs_m_thresholds_3_q0;
wire   [1:0] threshs_m_thresholds_2_address0;
reg    threshs_m_thresholds_2_ce0;
wire   [5:0] threshs_m_thresholds_2_q0;
wire   [1:0] threshs_m_thresholds_1_address0;
reg    threshs_m_thresholds_1_ce0;
wire   [5:0] threshs_m_thresholds_1_q0;
wire   [1:0] threshs_m_thresholds_address0;
reg    threshs_m_thresholds_ce0;
wire   [5:0] threshs_m_thresholds_q0;
wire   [1:0] threshs_m_thresholds_251_address0;
reg    threshs_m_thresholds_251_ce0;
wire   [5:0] threshs_m_thresholds_251_q0;
wire   [1:0] threshs_m_thresholds_250_address0;
reg    threshs_m_thresholds_250_ce0;
wire   [5:0] threshs_m_thresholds_250_q0;
wire   [1:0] threshs_m_thresholds_249_address0;
reg    threshs_m_thresholds_249_ce0;
wire   [5:0] threshs_m_thresholds_249_q0;
wire   [1:0] threshs_m_thresholds_248_address0;
reg    threshs_m_thresholds_248_ce0;
wire   [5:0] threshs_m_thresholds_248_q0;
wire   [1:0] threshs_m_thresholds_247_address0;
reg    threshs_m_thresholds_247_ce0;
wire   [5:0] threshs_m_thresholds_247_q0;
wire   [1:0] threshs_m_thresholds_246_address0;
reg    threshs_m_thresholds_246_ce0;
wire   [5:0] threshs_m_thresholds_246_q0;
wire   [1:0] threshs_m_thresholds_245_address0;
reg    threshs_m_thresholds_245_ce0;
wire   [5:0] threshs_m_thresholds_245_q0;
wire   [1:0] threshs_m_thresholds_244_address0;
reg    threshs_m_thresholds_244_ce0;
wire   [5:0] threshs_m_thresholds_244_q0;
wire   [1:0] threshs_m_thresholds_243_address0;
reg    threshs_m_thresholds_243_ce0;
wire   [5:0] threshs_m_thresholds_243_q0;
wire   [1:0] threshs_m_thresholds_242_address0;
reg    threshs_m_thresholds_242_ce0;
wire   [5:0] threshs_m_thresholds_242_q0;
wire   [1:0] threshs_m_thresholds_240_address0;
reg    threshs_m_thresholds_240_ce0;
wire   [5:0] threshs_m_thresholds_240_q0;
wire   [1:0] threshs_m_thresholds_239_address0;
reg    threshs_m_thresholds_239_ce0;
wire   [4:0] threshs_m_thresholds_239_q0;
wire   [1:0] threshs_m_thresholds_238_address0;
reg    threshs_m_thresholds_238_ce0;
wire   [4:0] threshs_m_thresholds_238_q0;
wire   [1:0] threshs_m_thresholds_237_address0;
reg    threshs_m_thresholds_237_ce0;
wire   [4:0] threshs_m_thresholds_237_q0;
wire   [1:0] threshs_m_thresholds_236_address0;
reg    threshs_m_thresholds_236_ce0;
wire   [4:0] threshs_m_thresholds_236_q0;
wire   [1:0] threshs_m_thresholds_235_address0;
reg    threshs_m_thresholds_235_ce0;
wire   [4:0] threshs_m_thresholds_235_q0;
wire   [1:0] threshs_m_thresholds_234_address0;
reg    threshs_m_thresholds_234_ce0;
wire   [4:0] threshs_m_thresholds_234_q0;
wire   [1:0] threshs_m_thresholds_233_address0;
reg    threshs_m_thresholds_233_ce0;
wire   [4:0] threshs_m_thresholds_233_q0;
wire   [1:0] threshs_m_thresholds_232_address0;
reg    threshs_m_thresholds_232_ce0;
wire   [4:0] threshs_m_thresholds_232_q0;
wire   [1:0] threshs_m_thresholds_231_address0;
reg    threshs_m_thresholds_231_ce0;
wire   [3:0] threshs_m_thresholds_231_q0;
wire   [1:0] threshs_m_thresholds_229_address0;
reg    threshs_m_thresholds_229_ce0;
wire   [3:0] threshs_m_thresholds_229_q0;
wire   [1:0] threshs_m_thresholds_228_address0;
reg    threshs_m_thresholds_228_ce0;
wire   [3:0] threshs_m_thresholds_228_q0;
wire   [1:0] threshs_m_thresholds_227_address0;
reg    threshs_m_thresholds_227_ce0;
wire   [3:0] threshs_m_thresholds_227_q0;
wire   [1:0] threshs_m_thresholds_226_address0;
reg    threshs_m_thresholds_226_ce0;
wire   [2:0] threshs_m_thresholds_226_q0;
wire   [1:0] threshs_m_thresholds_225_address0;
reg    threshs_m_thresholds_225_ce0;
wire   [2:0] threshs_m_thresholds_225_q0;
wire   [1:0] threshs_m_thresholds_224_address0;
reg    threshs_m_thresholds_224_ce0;
wire   [1:0] threshs_m_thresholds_224_q0;
wire   [1:0] threshs_m_thresholds_223_address0;
reg    threshs_m_thresholds_223_ce0;
wire   [0:0] threshs_m_thresholds_223_q0;
wire   [1:0] threshs_m_thresholds_222_address0;
reg    threshs_m_thresholds_222_ce0;
wire   [7:0] threshs_m_thresholds_222_q0;
wire   [1:0] threshs_m_thresholds_221_address0;
reg    threshs_m_thresholds_221_ce0;
wire   [7:0] threshs_m_thresholds_221_q0;
wire   [1:0] threshs_m_thresholds_220_address0;
reg    threshs_m_thresholds_220_ce0;
wire   [7:0] threshs_m_thresholds_220_q0;
wire   [1:0] threshs_m_thresholds_218_address0;
reg    threshs_m_thresholds_218_ce0;
wire   [7:0] threshs_m_thresholds_218_q0;
wire   [1:0] threshs_m_thresholds_217_address0;
reg    threshs_m_thresholds_217_ce0;
wire   [7:0] threshs_m_thresholds_217_q0;
wire   [1:0] threshs_m_thresholds_216_address0;
reg    threshs_m_thresholds_216_ce0;
wire   [7:0] threshs_m_thresholds_216_q0;
wire   [1:0] threshs_m_thresholds_215_address0;
reg    threshs_m_thresholds_215_ce0;
wire   [7:0] threshs_m_thresholds_215_q0;
wire   [1:0] threshs_m_thresholds_214_address0;
reg    threshs_m_thresholds_214_ce0;
wire   [7:0] threshs_m_thresholds_214_q0;
wire   [1:0] threshs_m_thresholds_213_address0;
reg    threshs_m_thresholds_213_ce0;
wire   [7:0] threshs_m_thresholds_213_q0;
wire   [1:0] threshs_m_thresholds_212_address0;
reg    threshs_m_thresholds_212_ce0;
wire   [7:0] threshs_m_thresholds_212_q0;
wire   [1:0] threshs_m_thresholds_211_address0;
reg    threshs_m_thresholds_211_ce0;
wire   [7:0] threshs_m_thresholds_211_q0;
wire   [1:0] threshs_m_thresholds_210_address0;
reg    threshs_m_thresholds_210_ce0;
wire   [7:0] threshs_m_thresholds_210_q0;
wire   [1:0] threshs_m_thresholds_209_address0;
reg    threshs_m_thresholds_209_ce0;
wire   [7:0] threshs_m_thresholds_209_q0;
wire   [1:0] threshs_m_thresholds_207_address0;
reg    threshs_m_thresholds_207_ce0;
wire   [7:0] threshs_m_thresholds_207_q0;
wire   [1:0] threshs_m_thresholds_206_address0;
reg    threshs_m_thresholds_206_ce0;
wire   [7:0] threshs_m_thresholds_206_q0;
wire   [1:0] threshs_m_thresholds_205_address0;
reg    threshs_m_thresholds_205_ce0;
wire   [7:0] threshs_m_thresholds_205_q0;
wire   [1:0] threshs_m_thresholds_204_address0;
reg    threshs_m_thresholds_204_ce0;
wire   [7:0] threshs_m_thresholds_204_q0;
wire   [1:0] threshs_m_thresholds_203_address0;
reg    threshs_m_thresholds_203_ce0;
wire   [7:0] threshs_m_thresholds_203_q0;
wire   [1:0] threshs_m_thresholds_202_address0;
reg    threshs_m_thresholds_202_ce0;
wire   [7:0] threshs_m_thresholds_202_q0;
wire   [1:0] threshs_m_thresholds_201_address0;
reg    threshs_m_thresholds_201_ce0;
wire   [7:0] threshs_m_thresholds_201_q0;
wire   [1:0] threshs_m_thresholds_200_address0;
reg    threshs_m_thresholds_200_ce0;
wire   [7:0] threshs_m_thresholds_200_q0;
wire   [1:0] threshs_m_thresholds_199_address0;
reg    threshs_m_thresholds_199_ce0;
wire   [7:0] threshs_m_thresholds_199_q0;
wire   [1:0] threshs_m_thresholds_198_address0;
reg    threshs_m_thresholds_198_ce0;
wire   [7:0] threshs_m_thresholds_198_q0;
wire   [1:0] threshs_m_thresholds_196_address0;
reg    threshs_m_thresholds_196_ce0;
wire   [7:0] threshs_m_thresholds_196_q0;
wire   [1:0] threshs_m_thresholds_195_address0;
reg    threshs_m_thresholds_195_ce0;
wire   [7:0] threshs_m_thresholds_195_q0;
wire   [1:0] threshs_m_thresholds_194_address0;
reg    threshs_m_thresholds_194_ce0;
wire   [7:0] threshs_m_thresholds_194_q0;
wire   [1:0] threshs_m_thresholds_193_address0;
reg    threshs_m_thresholds_193_ce0;
wire   [7:0] threshs_m_thresholds_193_q0;
wire   [1:0] threshs_m_thresholds_192_address0;
reg    threshs_m_thresholds_192_ce0;
wire   [7:0] threshs_m_thresholds_192_q0;
wire   [1:0] threshs_m_thresholds_191_address0;
reg    threshs_m_thresholds_191_ce0;
wire   [7:0] threshs_m_thresholds_191_q0;
wire   [1:0] threshs_m_thresholds_190_address0;
reg    threshs_m_thresholds_190_ce0;
wire   [7:0] threshs_m_thresholds_190_q0;
wire   [1:0] threshs_m_thresholds_189_address0;
reg    threshs_m_thresholds_189_ce0;
wire   [7:0] threshs_m_thresholds_189_q0;
wire   [1:0] threshs_m_thresholds_188_address0;
reg    threshs_m_thresholds_188_ce0;
wire   [7:0] threshs_m_thresholds_188_q0;
wire   [1:0] threshs_m_thresholds_187_address0;
reg    threshs_m_thresholds_187_ce0;
wire   [7:0] threshs_m_thresholds_187_q0;
wire   [1:0] threshs_m_thresholds_185_address0;
reg    threshs_m_thresholds_185_ce0;
wire   [7:0] threshs_m_thresholds_185_q0;
wire   [1:0] threshs_m_thresholds_184_address0;
reg    threshs_m_thresholds_184_ce0;
wire   [7:0] threshs_m_thresholds_184_q0;
wire   [1:0] threshs_m_thresholds_183_address0;
reg    threshs_m_thresholds_183_ce0;
wire   [7:0] threshs_m_thresholds_183_q0;
wire   [1:0] threshs_m_thresholds_182_address0;
reg    threshs_m_thresholds_182_ce0;
wire   [7:0] threshs_m_thresholds_182_q0;
wire   [1:0] threshs_m_thresholds_181_address0;
reg    threshs_m_thresholds_181_ce0;
wire   [7:0] threshs_m_thresholds_181_q0;
wire   [1:0] threshs_m_thresholds_180_address0;
reg    threshs_m_thresholds_180_ce0;
wire   [7:0] threshs_m_thresholds_180_q0;
wire   [1:0] threshs_m_thresholds_179_address0;
reg    threshs_m_thresholds_179_ce0;
wire   [7:0] threshs_m_thresholds_179_q0;
wire   [1:0] threshs_m_thresholds_178_address0;
reg    threshs_m_thresholds_178_ce0;
wire   [7:0] threshs_m_thresholds_178_q0;
wire   [1:0] threshs_m_thresholds_177_address0;
reg    threshs_m_thresholds_177_ce0;
wire   [7:0] threshs_m_thresholds_177_q0;
wire   [1:0] threshs_m_thresholds_176_address0;
reg    threshs_m_thresholds_176_ce0;
wire   [7:0] threshs_m_thresholds_176_q0;
wire   [1:0] threshs_m_thresholds_174_address0;
reg    threshs_m_thresholds_174_ce0;
wire   [7:0] threshs_m_thresholds_174_q0;
wire   [1:0] threshs_m_thresholds_173_address0;
reg    threshs_m_thresholds_173_ce0;
wire   [7:0] threshs_m_thresholds_173_q0;
wire   [1:0] threshs_m_thresholds_172_address0;
reg    threshs_m_thresholds_172_ce0;
wire   [7:0] threshs_m_thresholds_172_q0;
wire   [1:0] threshs_m_thresholds_171_address0;
reg    threshs_m_thresholds_171_ce0;
wire   [7:0] threshs_m_thresholds_171_q0;
wire   [1:0] threshs_m_thresholds_170_address0;
reg    threshs_m_thresholds_170_ce0;
wire   [7:0] threshs_m_thresholds_170_q0;
wire   [1:0] threshs_m_thresholds_169_address0;
reg    threshs_m_thresholds_169_ce0;
wire   [7:0] threshs_m_thresholds_169_q0;
wire   [1:0] threshs_m_thresholds_168_address0;
reg    threshs_m_thresholds_168_ce0;
wire   [7:0] threshs_m_thresholds_168_q0;
wire   [1:0] threshs_m_thresholds_167_address0;
reg    threshs_m_thresholds_167_ce0;
wire   [7:0] threshs_m_thresholds_167_q0;
wire   [1:0] threshs_m_thresholds_166_address0;
reg    threshs_m_thresholds_166_ce0;
wire   [7:0] threshs_m_thresholds_166_q0;
wire   [1:0] threshs_m_thresholds_165_address0;
reg    threshs_m_thresholds_165_ce0;
wire   [7:0] threshs_m_thresholds_165_q0;
wire   [1:0] threshs_m_thresholds_163_address0;
reg    threshs_m_thresholds_163_ce0;
wire   [7:0] threshs_m_thresholds_163_q0;
wire   [1:0] threshs_m_thresholds_162_address0;
reg    threshs_m_thresholds_162_ce0;
wire   [7:0] threshs_m_thresholds_162_q0;
wire   [1:0] threshs_m_thresholds_161_address0;
reg    threshs_m_thresholds_161_ce0;
wire   [7:0] threshs_m_thresholds_161_q0;
wire   [1:0] threshs_m_thresholds_160_address0;
reg    threshs_m_thresholds_160_ce0;
wire   [7:0] threshs_m_thresholds_160_q0;
wire   [1:0] threshs_m_thresholds_159_address0;
reg    threshs_m_thresholds_159_ce0;
wire   [7:0] threshs_m_thresholds_159_q0;
wire   [1:0] threshs_m_thresholds_158_address0;
reg    threshs_m_thresholds_158_ce0;
wire   [7:0] threshs_m_thresholds_158_q0;
wire   [1:0] threshs_m_thresholds_157_address0;
reg    threshs_m_thresholds_157_ce0;
wire   [7:0] threshs_m_thresholds_157_q0;
wire   [1:0] threshs_m_thresholds_156_address0;
reg    threshs_m_thresholds_156_ce0;
wire   [7:0] threshs_m_thresholds_156_q0;
wire   [1:0] threshs_m_thresholds_155_address0;
reg    threshs_m_thresholds_155_ce0;
wire   [7:0] threshs_m_thresholds_155_q0;
wire   [1:0] threshs_m_thresholds_154_address0;
reg    threshs_m_thresholds_154_ce0;
wire   [7:0] threshs_m_thresholds_154_q0;
wire   [1:0] threshs_m_thresholds_152_address0;
reg    threshs_m_thresholds_152_ce0;
wire   [7:0] threshs_m_thresholds_152_q0;
wire   [1:0] threshs_m_thresholds_151_address0;
reg    threshs_m_thresholds_151_ce0;
wire   [7:0] threshs_m_thresholds_151_q0;
wire   [1:0] threshs_m_thresholds_150_address0;
reg    threshs_m_thresholds_150_ce0;
wire   [6:0] threshs_m_thresholds_150_q0;
wire   [1:0] threshs_m_thresholds_149_address0;
reg    threshs_m_thresholds_149_ce0;
wire   [6:0] threshs_m_thresholds_149_q0;
wire   [1:0] threshs_m_thresholds_148_address0;
reg    threshs_m_thresholds_148_ce0;
wire   [6:0] threshs_m_thresholds_148_q0;
wire   [1:0] threshs_m_thresholds_147_address0;
reg    threshs_m_thresholds_147_ce0;
wire   [6:0] threshs_m_thresholds_147_q0;
wire   [1:0] threshs_m_thresholds_146_address0;
reg    threshs_m_thresholds_146_ce0;
wire   [6:0] threshs_m_thresholds_146_q0;
wire   [1:0] threshs_m_thresholds_145_address0;
reg    threshs_m_thresholds_145_ce0;
wire   [6:0] threshs_m_thresholds_145_q0;
wire   [1:0] threshs_m_thresholds_144_address0;
reg    threshs_m_thresholds_144_ce0;
wire   [6:0] threshs_m_thresholds_144_q0;
wire   [1:0] threshs_m_thresholds_143_address0;
reg    threshs_m_thresholds_143_ce0;
wire   [6:0] threshs_m_thresholds_143_q0;
wire   [1:0] threshs_m_thresholds_140_address0;
reg    threshs_m_thresholds_140_ce0;
wire   [6:0] threshs_m_thresholds_140_q0;
wire   [1:0] threshs_m_thresholds_139_address0;
reg    threshs_m_thresholds_139_ce0;
wire   [6:0] threshs_m_thresholds_139_q0;
wire   [1:0] threshs_m_thresholds_138_address0;
reg    threshs_m_thresholds_138_ce0;
wire   [6:0] threshs_m_thresholds_138_q0;
wire   [1:0] threshs_m_thresholds_137_address0;
reg    threshs_m_thresholds_137_ce0;
wire   [6:0] threshs_m_thresholds_137_q0;
wire   [1:0] threshs_m_thresholds_136_address0;
reg    threshs_m_thresholds_136_ce0;
wire   [6:0] threshs_m_thresholds_136_q0;
wire   [1:0] threshs_m_thresholds_135_address0;
reg    threshs_m_thresholds_135_ce0;
wire   [6:0] threshs_m_thresholds_135_q0;
wire   [1:0] threshs_m_thresholds_134_address0;
reg    threshs_m_thresholds_134_ce0;
wire   [6:0] threshs_m_thresholds_134_q0;
wire   [1:0] threshs_m_thresholds_133_address0;
reg    threshs_m_thresholds_133_ce0;
wire   [6:0] threshs_m_thresholds_133_q0;
wire   [1:0] threshs_m_thresholds_132_address0;
reg    threshs_m_thresholds_132_ce0;
wire   [6:0] threshs_m_thresholds_132_q0;
wire   [1:0] threshs_m_thresholds_131_address0;
reg    threshs_m_thresholds_131_ce0;
wire   [6:0] threshs_m_thresholds_131_q0;
wire   [1:0] threshs_m_thresholds_129_address0;
reg    threshs_m_thresholds_129_ce0;
wire   [6:0] threshs_m_thresholds_129_q0;
wire   [1:0] threshs_m_thresholds_128_address0;
reg    threshs_m_thresholds_128_ce0;
wire   [6:0] threshs_m_thresholds_128_q0;
wire   [1:0] threshs_m_thresholds_127_address0;
reg    threshs_m_thresholds_127_ce0;
wire   [6:0] threshs_m_thresholds_127_q0;
wire   [1:0] threshs_m_thresholds_126_address0;
reg    threshs_m_thresholds_126_ce0;
wire   [6:0] threshs_m_thresholds_126_q0;
wire   [1:0] threshs_m_thresholds_125_address0;
reg    threshs_m_thresholds_125_ce0;
wire   [6:0] threshs_m_thresholds_125_q0;
wire   [1:0] threshs_m_thresholds_124_address0;
reg    threshs_m_thresholds_124_ce0;
wire   [6:0] threshs_m_thresholds_124_q0;
wire   [1:0] threshs_m_thresholds_123_address0;
reg    threshs_m_thresholds_123_ce0;
wire   [6:0] threshs_m_thresholds_123_q0;
wire   [1:0] threshs_m_thresholds_122_address0;
reg    threshs_m_thresholds_122_ce0;
wire   [6:0] threshs_m_thresholds_122_q0;
wire   [1:0] threshs_m_thresholds_121_address0;
reg    threshs_m_thresholds_121_ce0;
wire   [6:0] threshs_m_thresholds_121_q0;
wire   [1:0] threshs_m_thresholds_120_address0;
reg    threshs_m_thresholds_120_ce0;
wire   [6:0] threshs_m_thresholds_120_q0;
wire   [1:0] threshs_m_thresholds_118_address0;
reg    threshs_m_thresholds_118_ce0;
wire   [6:0] threshs_m_thresholds_118_q0;
wire   [1:0] threshs_m_thresholds_117_address0;
reg    threshs_m_thresholds_117_ce0;
wire   [6:0] threshs_m_thresholds_117_q0;
wire   [1:0] threshs_m_thresholds_116_address0;
reg    threshs_m_thresholds_116_ce0;
wire   [6:0] threshs_m_thresholds_116_q0;
wire   [1:0] threshs_m_thresholds_115_address0;
reg    threshs_m_thresholds_115_ce0;
wire   [6:0] threshs_m_thresholds_115_q0;
wire   [1:0] threshs_m_thresholds_114_address0;
reg    threshs_m_thresholds_114_ce0;
wire   [5:0] threshs_m_thresholds_114_q0;
wire   [1:0] threshs_m_thresholds_113_address0;
reg    threshs_m_thresholds_113_ce0;
wire   [5:0] threshs_m_thresholds_113_q0;
wire   [1:0] threshs_m_thresholds_112_address0;
reg    threshs_m_thresholds_112_ce0;
wire   [5:0] threshs_m_thresholds_112_q0;
wire   [1:0] threshs_m_thresholds_111_address0;
reg    threshs_m_thresholds_111_ce0;
wire   [5:0] threshs_m_thresholds_111_q0;
wire   [1:0] threshs_m_thresholds_110_address0;
reg    threshs_m_thresholds_110_ce0;
wire   [5:0] threshs_m_thresholds_110_q0;
wire   [1:0] threshs_m_thresholds_109_address0;
reg    threshs_m_thresholds_109_ce0;
wire   [5:0] threshs_m_thresholds_109_q0;
wire   [1:0] threshs_m_thresholds_107_address0;
reg    threshs_m_thresholds_107_ce0;
wire   [5:0] threshs_m_thresholds_107_q0;
wire   [1:0] threshs_m_thresholds_106_address0;
reg    threshs_m_thresholds_106_ce0;
wire   [5:0] threshs_m_thresholds_106_q0;
wire   [1:0] threshs_m_thresholds_105_address0;
reg    threshs_m_thresholds_105_ce0;
wire   [5:0] threshs_m_thresholds_105_q0;
wire   [1:0] threshs_m_thresholds_104_address0;
reg    threshs_m_thresholds_104_ce0;
wire   [5:0] threshs_m_thresholds_104_q0;
wire   [1:0] threshs_m_thresholds_103_address0;
reg    threshs_m_thresholds_103_ce0;
wire   [5:0] threshs_m_thresholds_103_q0;
wire   [1:0] threshs_m_thresholds_102_address0;
reg    threshs_m_thresholds_102_ce0;
wire   [5:0] threshs_m_thresholds_102_q0;
wire   [1:0] threshs_m_thresholds_101_address0;
reg    threshs_m_thresholds_101_ce0;
wire   [5:0] threshs_m_thresholds_101_q0;
wire   [1:0] threshs_m_thresholds_100_address0;
reg    threshs_m_thresholds_100_ce0;
wire   [5:0] threshs_m_thresholds_100_q0;
wire   [1:0] threshs_m_thresholds_99_address0;
reg    threshs_m_thresholds_99_ce0;
wire   [5:0] threshs_m_thresholds_99_q0;
wire   [1:0] threshs_m_thresholds_98_address0;
reg    threshs_m_thresholds_98_ce0;
wire   [5:0] threshs_m_thresholds_98_q0;
wire   [1:0] threshs_m_thresholds_96_address0;
reg    threshs_m_thresholds_96_ce0;
wire   [4:0] threshs_m_thresholds_96_q0;
wire   [1:0] threshs_m_thresholds_95_address0;
reg    threshs_m_thresholds_95_ce0;
wire   [4:0] threshs_m_thresholds_95_q0;
wire   [1:0] threshs_m_thresholds_94_address0;
reg    threshs_m_thresholds_94_ce0;
wire   [4:0] threshs_m_thresholds_94_q0;
wire   [1:0] threshs_m_thresholds_93_address0;
reg    threshs_m_thresholds_93_ce0;
wire   [4:0] threshs_m_thresholds_93_q0;
wire   [1:0] threshs_m_thresholds_92_address0;
reg    threshs_m_thresholds_92_ce0;
wire   [4:0] threshs_m_thresholds_92_q0;
wire   [1:0] threshs_m_thresholds_91_address0;
reg    threshs_m_thresholds_91_ce0;
wire   [4:0] threshs_m_thresholds_91_q0;
wire   [1:0] threshs_m_thresholds_90_address0;
reg    threshs_m_thresholds_90_ce0;
wire   [4:0] threshs_m_thresholds_90_q0;
wire   [1:0] threshs_m_thresholds_89_address0;
reg    threshs_m_thresholds_89_ce0;
wire   [4:0] threshs_m_thresholds_89_q0;
wire   [1:0] threshs_m_thresholds_88_address0;
reg    threshs_m_thresholds_88_ce0;
wire   [3:0] threshs_m_thresholds_88_q0;
wire   [1:0] threshs_m_thresholds_87_address0;
reg    threshs_m_thresholds_87_ce0;
wire   [3:0] threshs_m_thresholds_87_q0;
wire   [1:0] threshs_m_thresholds_85_address0;
reg    threshs_m_thresholds_85_ce0;
wire   [3:0] threshs_m_thresholds_85_q0;
wire   [1:0] threshs_m_thresholds_84_address0;
reg    threshs_m_thresholds_84_ce0;
wire   [3:0] threshs_m_thresholds_84_q0;
wire   [1:0] threshs_m_thresholds_83_address0;
reg    threshs_m_thresholds_83_ce0;
wire   [2:0] threshs_m_thresholds_83_q0;
wire   [1:0] threshs_m_thresholds_82_address0;
reg    threshs_m_thresholds_82_ce0;
wire   [2:0] threshs_m_thresholds_82_q0;
wire   [1:0] threshs_m_thresholds_81_address0;
reg    threshs_m_thresholds_81_ce0;
wire   [1:0] threshs_m_thresholds_81_q0;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln221_fu_3928_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter3;
reg   [0:0] icmp_ln221_reg_11497;
reg   [0:0] icmp_ln221_reg_11497_pp0_iter2_reg;
reg   [31:0] nf_assign_reg_3906;
reg   [11:0] i_0_reg_3917;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
reg    ap_block_state5_io;
reg    ap_block_pp0_stage0_11001;
reg   [0:0] icmp_ln221_reg_11497_pp0_iter1_reg;
wire   [11:0] i_fu_3934_p2;
reg   [7:0] tmp_V_1_reg_11506;
wire   [31:0] nf_1_fu_4211_p3;
wire   [0:0] icmp_ln899_fu_4223_p2;
reg   [0:0] icmp_ln899_reg_13045;
wire   [0:0] icmp_ln899_1_fu_4232_p2;
reg   [0:0] icmp_ln899_1_reg_13050;
wire   [0:0] icmp_ln899_2_fu_4245_p2;
reg   [0:0] icmp_ln899_2_reg_13055;
wire   [2:0] add_ln700_4_fu_9046_p2;
reg   [2:0] add_ln700_4_reg_13060;
wire   [2:0] add_ln700_8_fu_9072_p2;
reg   [2:0] add_ln700_8_reg_13065;
wire   [2:0] add_ln700_11_fu_9098_p2;
reg   [2:0] add_ln700_11_reg_13070;
wire   [2:0] add_ln700_16_fu_9124_p2;
reg   [2:0] add_ln700_16_reg_13075;
wire   [2:0] add_ln700_19_fu_9150_p2;
reg   [2:0] add_ln700_19_reg_13080;
wire   [2:0] add_ln700_23_fu_9176_p2;
reg   [2:0] add_ln700_23_reg_13085;
wire   [2:0] add_ln700_26_fu_9202_p2;
reg   [2:0] add_ln700_26_reg_13090;
wire   [2:0] add_ln700_32_fu_9228_p2;
reg   [2:0] add_ln700_32_reg_13095;
wire   [2:0] add_ln700_35_fu_9254_p2;
reg   [2:0] add_ln700_35_reg_13100;
wire   [2:0] add_ln700_39_fu_9280_p2;
reg   [2:0] add_ln700_39_reg_13105;
wire   [2:0] add_ln700_42_fu_9306_p2;
reg   [2:0] add_ln700_42_reg_13110;
wire   [2:0] add_ln700_47_fu_9332_p2;
reg   [2:0] add_ln700_47_reg_13115;
wire   [2:0] add_ln700_50_fu_9358_p2;
reg   [2:0] add_ln700_50_reg_13120;
wire   [2:0] add_ln700_54_fu_9384_p2;
reg   [2:0] add_ln700_54_reg_13125;
wire   [2:0] add_ln700_57_fu_9410_p2;
reg   [2:0] add_ln700_57_reg_13130;
wire   [2:0] add_ln700_64_fu_9436_p2;
reg   [2:0] add_ln700_64_reg_13135;
wire   [2:0] add_ln700_67_fu_9462_p2;
reg   [2:0] add_ln700_67_reg_13140;
wire   [2:0] add_ln700_71_fu_9488_p2;
reg   [2:0] add_ln700_71_reg_13145;
wire   [2:0] add_ln700_74_fu_9514_p2;
reg   [2:0] add_ln700_74_reg_13150;
wire   [2:0] add_ln700_79_fu_9540_p2;
reg   [2:0] add_ln700_79_reg_13155;
wire   [2:0] add_ln700_82_fu_9566_p2;
reg   [2:0] add_ln700_82_reg_13160;
wire   [2:0] add_ln700_86_fu_9592_p2;
reg   [2:0] add_ln700_86_reg_13165;
wire   [2:0] add_ln700_89_fu_9618_p2;
reg   [2:0] add_ln700_89_reg_13170;
wire   [2:0] add_ln700_95_fu_9644_p2;
reg   [2:0] add_ln700_95_reg_13175;
wire   [2:0] add_ln700_98_fu_9670_p2;
reg   [2:0] add_ln700_98_reg_13180;
wire   [2:0] add_ln700_102_fu_9696_p2;
reg   [2:0] add_ln700_102_reg_13185;
wire   [2:0] add_ln700_105_fu_9722_p2;
reg   [2:0] add_ln700_105_reg_13190;
wire   [2:0] add_ln700_110_fu_9748_p2;
reg   [2:0] add_ln700_110_reg_13195;
wire   [2:0] add_ln700_113_fu_9774_p2;
reg   [2:0] add_ln700_113_reg_13200;
wire   [2:0] add_ln700_117_fu_9800_p2;
reg   [2:0] add_ln700_117_reg_13205;
wire   [2:0] add_ln700_120_fu_9826_p2;
reg   [2:0] add_ln700_120_reg_13210;
wire   [2:0] add_ln700_128_fu_9852_p2;
reg   [2:0] add_ln700_128_reg_13215;
wire   [2:0] add_ln700_131_fu_9878_p2;
reg   [2:0] add_ln700_131_reg_13220;
wire   [2:0] add_ln700_135_fu_9904_p2;
reg   [2:0] add_ln700_135_reg_13225;
wire   [2:0] add_ln700_138_fu_9930_p2;
reg   [2:0] add_ln700_138_reg_13230;
wire   [2:0] add_ln700_143_fu_9956_p2;
reg   [2:0] add_ln700_143_reg_13235;
wire   [2:0] add_ln700_146_fu_9982_p2;
reg   [2:0] add_ln700_146_reg_13240;
wire   [2:0] add_ln700_150_fu_10008_p2;
reg   [2:0] add_ln700_150_reg_13245;
wire   [2:0] add_ln700_153_fu_10034_p2;
reg   [2:0] add_ln700_153_reg_13250;
wire   [2:0] add_ln700_159_fu_10060_p2;
reg   [2:0] add_ln700_159_reg_13255;
wire   [2:0] add_ln700_162_fu_10086_p2;
reg   [2:0] add_ln700_162_reg_13260;
wire   [2:0] add_ln700_166_fu_10112_p2;
reg   [2:0] add_ln700_166_reg_13265;
wire   [2:0] add_ln700_169_fu_10138_p2;
reg   [2:0] add_ln700_169_reg_13270;
wire   [2:0] add_ln700_174_fu_10164_p2;
reg   [2:0] add_ln700_174_reg_13275;
wire   [2:0] add_ln700_177_fu_10190_p2;
reg   [2:0] add_ln700_177_reg_13280;
wire   [2:0] add_ln700_181_fu_10216_p2;
reg   [2:0] add_ln700_181_reg_13285;
wire   [2:0] add_ln700_184_fu_10242_p2;
reg   [2:0] add_ln700_184_reg_13290;
wire   [2:0] add_ln700_191_fu_10268_p2;
reg   [2:0] add_ln700_191_reg_13295;
wire   [2:0] add_ln700_194_fu_10294_p2;
reg   [2:0] add_ln700_194_reg_13300;
wire   [2:0] add_ln700_198_fu_10320_p2;
reg   [2:0] add_ln700_198_reg_13305;
wire   [2:0] add_ln700_201_fu_10346_p2;
reg   [2:0] add_ln700_201_reg_13310;
wire   [2:0] add_ln700_206_fu_10372_p2;
reg   [2:0] add_ln700_206_reg_13315;
wire   [2:0] add_ln700_209_fu_10398_p2;
reg   [2:0] add_ln700_209_reg_13320;
wire   [2:0] add_ln700_213_fu_10424_p2;
reg   [2:0] add_ln700_213_reg_13325;
wire   [2:0] add_ln700_216_fu_10450_p2;
reg   [2:0] add_ln700_216_reg_13330;
wire   [2:0] add_ln700_222_fu_10476_p2;
reg   [2:0] add_ln700_222_reg_13335;
wire   [2:0] add_ln700_225_fu_10502_p2;
reg   [2:0] add_ln700_225_reg_13340;
wire   [2:0] add_ln700_229_fu_10528_p2;
reg   [2:0] add_ln700_229_reg_13345;
wire   [2:0] add_ln700_232_fu_10554_p2;
reg   [2:0] add_ln700_232_reg_13350;
wire   [2:0] add_ln700_237_fu_10580_p2;
reg   [2:0] add_ln700_237_reg_13355;
wire   [2:0] add_ln700_240_fu_10606_p2;
reg   [2:0] add_ln700_240_reg_13360;
wire   [2:0] add_ln700_244_fu_10632_p2;
reg   [2:0] add_ln700_244_reg_13365;
wire   [2:0] add_ln700_247_fu_10658_p2;
reg   [2:0] add_ln700_247_reg_13370;
wire   [7:0] add_ln700_13_fu_10736_p2;
reg   [7:0] add_ln700_13_reg_13375;
wire   [4:0] add_ln700_28_fu_10774_p2;
reg   [4:0] add_ln700_28_reg_13380;
wire   [5:0] add_ln700_60_fu_10864_p2;
reg   [5:0] add_ln700_60_reg_13385;
wire   [6:0] add_ln700_124_fu_11058_p2;
reg   [6:0] add_ln700_124_reg_13390;
wire   [6:0] add_ln700_188_fu_11252_p2;
reg   [6:0] add_ln700_188_reg_13395;
wire   [6:0] add_ln700_251_fu_11446_p2;
reg   [6:0] add_ln700_251_reg_13400;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
wire   [63:0] zext_ln142_fu_3940_p1;
reg    ap_block_pp0_stage0_01001;
wire   [31:0] nf_fu_4199_p2;
wire   [0:0] icmp_ln235_fu_4205_p2;
wire   [7:0] zext_ln142_1_fu_4219_p1;
wire   [7:0] zext_ln142_2_fu_4228_p1;
wire   [7:0] select_ln142_fu_4237_p3;
wire   [7:0] zext_ln142_5_fu_4250_p1;
wire   [0:0] icmp_ln899_3_fu_4254_p2;
wire   [0:0] xor_ln899_3_fu_4259_p2;
wire   [7:0] zext_ln142_7_fu_4269_p1;
wire   [0:0] icmp_ln899_4_fu_4273_p2;
wire   [0:0] xor_ln899_4_fu_4278_p2;
wire  signed [2:0] sext_ln142_fu_4288_p1;
wire   [7:0] zext_ln142_9_fu_4292_p1;
wire   [0:0] icmp_ln899_5_fu_4296_p2;
wire   [0:0] xor_ln899_5_fu_4301_p2;
wire   [7:0] select_ln142_1_fu_4311_p3;
wire   [0:0] icmp_ln899_6_fu_4319_p2;
wire   [0:0] xor_ln899_6_fu_4324_p2;
wire   [7:0] zext_ln142_12_fu_4334_p1;
wire   [0:0] icmp_ln899_7_fu_4338_p2;
wire   [0:0] xor_ln899_7_fu_4343_p2;
wire   [7:0] zext_ln142_14_fu_4353_p1;
wire   [0:0] icmp_ln899_8_fu_4357_p2;
wire   [0:0] xor_ln899_8_fu_4362_p2;
wire   [7:0] zext_ln142_16_fu_4372_p1;
wire   [0:0] icmp_ln899_9_fu_4376_p2;
wire   [0:0] xor_ln899_9_fu_4381_p2;
wire   [7:0] zext_ln142_18_fu_4391_p1;
wire   [0:0] icmp_ln899_10_fu_4395_p2;
wire   [0:0] xor_ln899_10_fu_4400_p2;
wire  signed [3:0] sext_ln142_1_fu_4410_p1;
wire   [7:0] zext_ln142_20_fu_4414_p1;
wire   [0:0] icmp_ln899_11_fu_4418_p2;
wire   [0:0] xor_ln899_11_fu_4423_p2;
wire  signed [3:0] sext_ln142_2_fu_4433_p1;
wire   [7:0] zext_ln142_22_fu_4437_p1;
wire   [0:0] icmp_ln899_12_fu_4441_p2;
wire   [0:0] xor_ln899_12_fu_4446_p2;
wire  signed [3:0] sext_ln142_3_fu_4456_p1;
wire   [7:0] zext_ln142_24_fu_4460_p1;
wire   [0:0] icmp_ln899_13_fu_4464_p2;
wire   [0:0] xor_ln899_13_fu_4469_p2;
wire   [7:0] select_ln142_2_fu_4479_p3;
wire   [0:0] icmp_ln899_14_fu_4487_p2;
wire   [0:0] xor_ln899_14_fu_4492_p2;
wire   [7:0] zext_ln142_27_fu_4502_p1;
wire   [0:0] icmp_ln899_15_fu_4506_p2;
wire   [0:0] xor_ln899_15_fu_4511_p2;
wire   [7:0] zext_ln142_29_fu_4521_p1;
wire   [0:0] icmp_ln899_16_fu_4525_p2;
wire   [0:0] xor_ln899_16_fu_4530_p2;
wire   [7:0] zext_ln142_31_fu_4540_p1;
wire   [0:0] icmp_ln899_17_fu_4544_p2;
wire   [0:0] xor_ln899_17_fu_4549_p2;
wire   [7:0] zext_ln142_33_fu_4559_p1;
wire   [0:0] icmp_ln899_18_fu_4563_p2;
wire   [0:0] xor_ln899_18_fu_4568_p2;
wire   [7:0] zext_ln142_35_fu_4578_p1;
wire   [0:0] icmp_ln899_19_fu_4582_p2;
wire   [0:0] xor_ln899_19_fu_4587_p2;
wire   [7:0] zext_ln142_37_fu_4597_p1;
wire   [0:0] icmp_ln899_20_fu_4601_p2;
wire   [0:0] xor_ln899_20_fu_4606_p2;
wire   [7:0] zext_ln142_39_fu_4616_p1;
wire   [0:0] icmp_ln899_21_fu_4620_p2;
wire   [0:0] xor_ln899_21_fu_4625_p2;
wire   [7:0] zext_ln142_41_fu_4635_p1;
wire   [0:0] icmp_ln899_22_fu_4639_p2;
wire   [0:0] xor_ln899_22_fu_4644_p2;
wire  signed [4:0] sext_ln142_4_fu_4654_p1;
wire   [7:0] zext_ln142_43_fu_4658_p1;
wire   [0:0] icmp_ln899_23_fu_4662_p2;
wire   [0:0] xor_ln899_23_fu_4667_p2;
wire  signed [4:0] sext_ln142_5_fu_4677_p1;
wire   [7:0] zext_ln142_45_fu_4681_p1;
wire   [0:0] icmp_ln899_24_fu_4685_p2;
wire   [0:0] xor_ln899_24_fu_4690_p2;
wire  signed [4:0] sext_ln142_6_fu_4700_p1;
wire   [7:0] zext_ln142_47_fu_4704_p1;
wire   [0:0] icmp_ln899_25_fu_4708_p2;
wire   [0:0] xor_ln899_25_fu_4713_p2;
wire  signed [4:0] sext_ln142_7_fu_4723_p1;
wire   [7:0] zext_ln142_49_fu_4727_p1;
wire   [0:0] icmp_ln899_26_fu_4731_p2;
wire   [0:0] xor_ln899_26_fu_4736_p2;
wire  signed [4:0] sext_ln142_8_fu_4746_p1;
wire   [7:0] zext_ln142_51_fu_4750_p1;
wire   [0:0] icmp_ln899_27_fu_4754_p2;
wire   [0:0] xor_ln899_27_fu_4759_p2;
wire  signed [4:0] sext_ln142_9_fu_4769_p1;
wire   [7:0] zext_ln142_53_fu_4773_p1;
wire   [0:0] icmp_ln899_28_fu_4777_p2;
wire   [0:0] xor_ln899_28_fu_4782_p2;
wire  signed [4:0] sext_ln142_10_fu_4792_p1;
wire   [7:0] zext_ln142_55_fu_4796_p1;
wire   [0:0] icmp_ln899_29_fu_4800_p2;
wire   [0:0] xor_ln899_29_fu_4805_p2;
wire   [7:0] select_ln142_3_fu_4815_p3;
wire   [0:0] icmp_ln899_30_fu_4823_p2;
wire   [0:0] xor_ln899_30_fu_4828_p2;
wire   [7:0] zext_ln142_58_fu_4838_p1;
wire   [0:0] icmp_ln899_31_fu_4842_p2;
wire   [0:0] xor_ln899_31_fu_4847_p2;
wire   [7:0] zext_ln142_60_fu_4857_p1;
wire   [0:0] icmp_ln899_32_fu_4861_p2;
wire   [0:0] xor_ln899_32_fu_4866_p2;
wire   [7:0] zext_ln142_62_fu_4876_p1;
wire   [0:0] icmp_ln899_33_fu_4880_p2;
wire   [0:0] xor_ln899_33_fu_4885_p2;
wire   [7:0] zext_ln142_64_fu_4895_p1;
wire   [0:0] icmp_ln899_34_fu_4899_p2;
wire   [0:0] xor_ln899_34_fu_4904_p2;
wire   [7:0] zext_ln142_66_fu_4914_p1;
wire   [0:0] icmp_ln899_35_fu_4918_p2;
wire   [0:0] xor_ln899_35_fu_4923_p2;
wire   [7:0] zext_ln142_68_fu_4933_p1;
wire   [0:0] icmp_ln899_36_fu_4937_p2;
wire   [0:0] xor_ln899_36_fu_4942_p2;
wire   [7:0] zext_ln142_70_fu_4952_p1;
wire   [0:0] icmp_ln899_37_fu_4956_p2;
wire   [0:0] xor_ln899_37_fu_4961_p2;
wire   [7:0] zext_ln142_72_fu_4971_p1;
wire   [0:0] icmp_ln899_38_fu_4975_p2;
wire   [0:0] xor_ln899_38_fu_4980_p2;
wire   [7:0] zext_ln142_74_fu_4990_p1;
wire   [0:0] icmp_ln899_39_fu_4994_p2;
wire   [0:0] xor_ln899_39_fu_4999_p2;
wire   [7:0] zext_ln142_76_fu_5009_p1;
wire   [0:0] icmp_ln899_40_fu_5013_p2;
wire   [0:0] xor_ln899_40_fu_5018_p2;
wire   [7:0] zext_ln142_78_fu_5028_p1;
wire   [0:0] icmp_ln899_41_fu_5032_p2;
wire   [0:0] xor_ln899_41_fu_5037_p2;
wire   [7:0] zext_ln142_80_fu_5047_p1;
wire   [0:0] icmp_ln899_42_fu_5051_p2;
wire   [0:0] xor_ln899_42_fu_5056_p2;
wire   [7:0] zext_ln142_82_fu_5066_p1;
wire   [0:0] icmp_ln899_43_fu_5070_p2;
wire   [0:0] xor_ln899_43_fu_5075_p2;
wire   [7:0] zext_ln142_84_fu_5085_p1;
wire   [0:0] icmp_ln899_44_fu_5089_p2;
wire   [0:0] xor_ln899_44_fu_5094_p2;
wire   [7:0] zext_ln142_86_fu_5104_p1;
wire   [0:0] icmp_ln899_45_fu_5108_p2;
wire   [0:0] xor_ln899_45_fu_5113_p2;
wire   [7:0] zext_ln142_88_fu_5123_p1;
wire   [0:0] icmp_ln899_46_fu_5127_p2;
wire   [0:0] xor_ln899_46_fu_5132_p2;
wire  signed [5:0] sext_ln142_11_fu_5142_p1;
wire   [7:0] zext_ln142_90_fu_5146_p1;
wire   [0:0] icmp_ln899_47_fu_5150_p2;
wire   [0:0] xor_ln899_47_fu_5155_p2;
wire  signed [5:0] sext_ln142_12_fu_5165_p1;
wire   [7:0] zext_ln142_92_fu_5169_p1;
wire   [0:0] icmp_ln899_48_fu_5173_p2;
wire   [0:0] xor_ln899_48_fu_5178_p2;
wire  signed [5:0] sext_ln142_13_fu_5188_p1;
wire   [7:0] zext_ln142_94_fu_5192_p1;
wire   [0:0] icmp_ln899_49_fu_5196_p2;
wire   [0:0] xor_ln899_49_fu_5201_p2;
wire  signed [5:0] sext_ln142_14_fu_5211_p1;
wire   [7:0] zext_ln142_96_fu_5215_p1;
wire   [0:0] icmp_ln899_50_fu_5219_p2;
wire   [0:0] xor_ln899_50_fu_5224_p2;
wire  signed [5:0] sext_ln142_15_fu_5234_p1;
wire   [7:0] zext_ln142_98_fu_5238_p1;
wire   [0:0] icmp_ln899_51_fu_5242_p2;
wire   [0:0] xor_ln899_51_fu_5247_p2;
wire  signed [5:0] sext_ln142_16_fu_5257_p1;
wire   [7:0] zext_ln142_100_fu_5261_p1;
wire   [0:0] icmp_ln899_52_fu_5265_p2;
wire   [0:0] xor_ln899_52_fu_5270_p2;
wire  signed [5:0] sext_ln142_17_fu_5280_p1;
wire   [7:0] zext_ln142_102_fu_5284_p1;
wire   [0:0] icmp_ln899_53_fu_5288_p2;
wire   [0:0] xor_ln899_53_fu_5293_p2;
wire  signed [5:0] sext_ln142_18_fu_5303_p1;
wire   [7:0] zext_ln142_104_fu_5307_p1;
wire   [0:0] icmp_ln899_54_fu_5311_p2;
wire   [0:0] xor_ln899_54_fu_5316_p2;
wire  signed [5:0] sext_ln142_19_fu_5326_p1;
wire   [7:0] zext_ln142_106_fu_5330_p1;
wire   [0:0] icmp_ln899_55_fu_5334_p2;
wire   [0:0] xor_ln899_55_fu_5339_p2;
wire  signed [5:0] sext_ln142_20_fu_5349_p1;
wire   [7:0] zext_ln142_108_fu_5353_p1;
wire   [0:0] icmp_ln899_56_fu_5357_p2;
wire   [0:0] xor_ln899_56_fu_5362_p2;
wire  signed [5:0] sext_ln142_21_fu_5372_p1;
wire   [7:0] zext_ln142_110_fu_5376_p1;
wire   [0:0] icmp_ln899_57_fu_5380_p2;
wire   [0:0] xor_ln899_57_fu_5385_p2;
wire  signed [5:0] sext_ln142_22_fu_5395_p1;
wire   [7:0] zext_ln142_112_fu_5399_p1;
wire   [0:0] icmp_ln899_58_fu_5403_p2;
wire   [0:0] xor_ln899_58_fu_5408_p2;
wire  signed [5:0] sext_ln142_23_fu_5418_p1;
wire   [7:0] zext_ln142_114_fu_5422_p1;
wire   [0:0] icmp_ln899_59_fu_5426_p2;
wire   [0:0] xor_ln899_59_fu_5431_p2;
wire  signed [5:0] sext_ln142_24_fu_5441_p1;
wire   [7:0] zext_ln142_116_fu_5445_p1;
wire   [0:0] icmp_ln899_60_fu_5449_p2;
wire   [0:0] xor_ln899_60_fu_5454_p2;
wire  signed [5:0] sext_ln142_25_fu_5464_p1;
wire   [7:0] zext_ln142_118_fu_5468_p1;
wire   [0:0] icmp_ln899_61_fu_5472_p2;
wire   [0:0] xor_ln899_61_fu_5477_p2;
wire   [7:0] select_ln142_4_fu_5487_p3;
wire   [0:0] icmp_ln899_62_fu_5495_p2;
wire   [0:0] xor_ln899_62_fu_5500_p2;
wire   [7:0] zext_ln142_121_fu_5510_p1;
wire   [0:0] icmp_ln899_63_fu_5514_p2;
wire   [0:0] xor_ln899_63_fu_5519_p2;
wire   [7:0] zext_ln142_123_fu_5529_p1;
wire   [0:0] icmp_ln899_64_fu_5533_p2;
wire   [0:0] xor_ln899_64_fu_5538_p2;
wire   [7:0] zext_ln142_125_fu_5548_p1;
wire   [0:0] icmp_ln899_65_fu_5552_p2;
wire   [0:0] xor_ln899_65_fu_5557_p2;
wire   [7:0] zext_ln142_127_fu_5567_p1;
wire   [0:0] icmp_ln899_66_fu_5571_p2;
wire   [0:0] xor_ln899_66_fu_5576_p2;
wire   [7:0] zext_ln142_129_fu_5586_p1;
wire   [0:0] icmp_ln899_67_fu_5590_p2;
wire   [0:0] xor_ln899_67_fu_5595_p2;
wire   [7:0] zext_ln142_131_fu_5605_p1;
wire   [0:0] icmp_ln899_68_fu_5609_p2;
wire   [0:0] xor_ln899_68_fu_5614_p2;
wire   [7:0] zext_ln142_133_fu_5624_p1;
wire   [0:0] icmp_ln899_69_fu_5628_p2;
wire   [0:0] xor_ln899_69_fu_5633_p2;
wire   [7:0] zext_ln142_135_fu_5643_p1;
wire   [0:0] icmp_ln899_70_fu_5647_p2;
wire   [0:0] xor_ln899_70_fu_5652_p2;
wire   [7:0] zext_ln142_137_fu_5662_p1;
wire   [0:0] icmp_ln899_71_fu_5666_p2;
wire   [0:0] xor_ln899_71_fu_5671_p2;
wire   [7:0] zext_ln142_139_fu_5681_p1;
wire   [0:0] icmp_ln899_72_fu_5685_p2;
wire   [0:0] xor_ln899_72_fu_5690_p2;
wire   [7:0] zext_ln142_141_fu_5700_p1;
wire   [0:0] icmp_ln899_73_fu_5704_p2;
wire   [0:0] xor_ln899_73_fu_5709_p2;
wire   [7:0] zext_ln142_143_fu_5719_p1;
wire   [0:0] icmp_ln899_74_fu_5723_p2;
wire   [0:0] xor_ln899_74_fu_5728_p2;
wire   [7:0] zext_ln142_145_fu_5738_p1;
wire   [0:0] icmp_ln899_75_fu_5742_p2;
wire   [0:0] xor_ln899_75_fu_5747_p2;
wire   [7:0] zext_ln142_147_fu_5757_p1;
wire   [0:0] icmp_ln899_76_fu_5761_p2;
wire   [0:0] xor_ln899_76_fu_5766_p2;
wire   [7:0] zext_ln142_149_fu_5776_p1;
wire   [0:0] icmp_ln899_77_fu_5780_p2;
wire   [0:0] xor_ln899_77_fu_5785_p2;
wire   [7:0] zext_ln142_151_fu_5795_p1;
wire   [0:0] icmp_ln899_78_fu_5799_p2;
wire   [0:0] xor_ln899_78_fu_5804_p2;
wire   [7:0] zext_ln142_153_fu_5814_p1;
wire   [0:0] icmp_ln899_79_fu_5818_p2;
wire   [0:0] xor_ln899_79_fu_5823_p2;
wire   [7:0] zext_ln142_155_fu_5833_p1;
wire   [0:0] icmp_ln899_80_fu_5837_p2;
wire   [0:0] xor_ln899_80_fu_5842_p2;
wire   [7:0] zext_ln142_157_fu_5852_p1;
wire   [0:0] icmp_ln899_81_fu_5856_p2;
wire   [0:0] xor_ln899_81_fu_5861_p2;
wire   [7:0] zext_ln142_159_fu_5871_p1;
wire   [0:0] icmp_ln899_82_fu_5875_p2;
wire   [0:0] xor_ln899_82_fu_5880_p2;
wire   [7:0] zext_ln142_161_fu_5890_p1;
wire   [0:0] icmp_ln899_83_fu_5894_p2;
wire   [0:0] xor_ln899_83_fu_5899_p2;
wire   [7:0] zext_ln142_163_fu_5909_p1;
wire   [0:0] icmp_ln899_84_fu_5913_p2;
wire   [0:0] xor_ln899_84_fu_5918_p2;
wire   [7:0] zext_ln142_165_fu_5928_p1;
wire   [0:0] icmp_ln899_85_fu_5932_p2;
wire   [0:0] xor_ln899_85_fu_5937_p2;
wire   [7:0] zext_ln142_167_fu_5947_p1;
wire   [0:0] icmp_ln899_86_fu_5951_p2;
wire   [0:0] xor_ln899_86_fu_5956_p2;
wire   [7:0] zext_ln142_169_fu_5966_p1;
wire   [0:0] icmp_ln899_87_fu_5970_p2;
wire   [0:0] xor_ln899_87_fu_5975_p2;
wire   [7:0] zext_ln142_171_fu_5985_p1;
wire   [0:0] icmp_ln899_88_fu_5989_p2;
wire   [0:0] xor_ln899_88_fu_5994_p2;
wire   [7:0] zext_ln142_173_fu_6004_p1;
wire   [0:0] icmp_ln899_89_fu_6008_p2;
wire   [0:0] xor_ln899_89_fu_6013_p2;
wire   [7:0] zext_ln142_175_fu_6023_p1;
wire   [0:0] icmp_ln899_90_fu_6027_p2;
wire   [0:0] xor_ln899_90_fu_6032_p2;
wire   [7:0] zext_ln142_177_fu_6042_p1;
wire   [0:0] icmp_ln899_91_fu_6046_p2;
wire   [0:0] xor_ln899_91_fu_6051_p2;
wire   [7:0] zext_ln142_179_fu_6061_p1;
wire   [0:0] icmp_ln899_92_fu_6065_p2;
wire   [0:0] xor_ln899_92_fu_6070_p2;
wire   [7:0] zext_ln142_181_fu_6080_p1;
wire   [0:0] icmp_ln899_93_fu_6084_p2;
wire   [0:0] xor_ln899_93_fu_6089_p2;
wire   [7:0] zext_ln142_183_fu_6099_p1;
wire   [0:0] icmp_ln899_94_fu_6103_p2;
wire   [0:0] xor_ln899_94_fu_6108_p2;
wire  signed [6:0] sext_ln142_26_fu_6118_p1;
wire   [7:0] zext_ln142_185_fu_6122_p1;
wire   [0:0] icmp_ln899_95_fu_6126_p2;
wire   [0:0] xor_ln899_95_fu_6131_p2;
wire  signed [6:0] sext_ln142_27_fu_6141_p1;
wire   [7:0] zext_ln142_187_fu_6145_p1;
wire   [0:0] icmp_ln899_96_fu_6149_p2;
wire   [0:0] xor_ln899_96_fu_6154_p2;
wire  signed [6:0] sext_ln142_28_fu_6164_p1;
wire   [7:0] zext_ln142_189_fu_6168_p1;
wire   [0:0] icmp_ln899_97_fu_6172_p2;
wire   [0:0] xor_ln899_97_fu_6177_p2;
wire  signed [6:0] sext_ln142_29_fu_6187_p1;
wire   [7:0] zext_ln142_191_fu_6191_p1;
wire   [0:0] icmp_ln899_98_fu_6195_p2;
wire   [0:0] xor_ln899_98_fu_6200_p2;
wire  signed [6:0] sext_ln142_30_fu_6210_p1;
wire   [7:0] zext_ln142_193_fu_6214_p1;
wire   [0:0] icmp_ln899_99_fu_6218_p2;
wire   [0:0] xor_ln899_99_fu_6223_p2;
wire  signed [6:0] sext_ln142_31_fu_6233_p1;
wire   [7:0] zext_ln142_195_fu_6237_p1;
wire   [0:0] icmp_ln899_100_fu_6241_p2;
wire   [0:0] xor_ln899_100_fu_6246_p2;
wire  signed [6:0] sext_ln142_32_fu_6256_p1;
wire   [7:0] zext_ln142_197_fu_6260_p1;
wire   [0:0] icmp_ln899_101_fu_6264_p2;
wire   [0:0] xor_ln899_101_fu_6269_p2;
wire  signed [6:0] sext_ln142_33_fu_6279_p1;
wire   [7:0] zext_ln142_199_fu_6283_p1;
wire   [0:0] icmp_ln899_102_fu_6287_p2;
wire   [0:0] xor_ln899_102_fu_6292_p2;
wire  signed [6:0] sext_ln142_34_fu_6302_p1;
wire   [7:0] zext_ln142_201_fu_6306_p1;
wire   [0:0] icmp_ln899_103_fu_6310_p2;
wire   [0:0] xor_ln899_103_fu_6315_p2;
wire  signed [6:0] sext_ln142_35_fu_6325_p1;
wire   [7:0] zext_ln142_203_fu_6329_p1;
wire   [0:0] icmp_ln899_104_fu_6333_p2;
wire   [0:0] xor_ln899_104_fu_6338_p2;
wire  signed [6:0] sext_ln142_36_fu_6348_p1;
wire   [7:0] zext_ln142_205_fu_6352_p1;
wire   [0:0] icmp_ln899_105_fu_6356_p2;
wire   [0:0] xor_ln899_105_fu_6361_p2;
wire  signed [6:0] sext_ln142_37_fu_6371_p1;
wire   [7:0] zext_ln142_207_fu_6375_p1;
wire   [0:0] icmp_ln899_106_fu_6379_p2;
wire   [0:0] xor_ln899_106_fu_6384_p2;
wire  signed [6:0] sext_ln142_38_fu_6394_p1;
wire   [7:0] zext_ln142_209_fu_6398_p1;
wire   [0:0] icmp_ln899_107_fu_6402_p2;
wire   [0:0] xor_ln899_107_fu_6407_p2;
wire  signed [6:0] sext_ln142_39_fu_6417_p1;
wire   [7:0] zext_ln142_211_fu_6421_p1;
wire   [0:0] icmp_ln899_108_fu_6425_p2;
wire   [0:0] xor_ln899_108_fu_6430_p2;
wire  signed [6:0] sext_ln142_40_fu_6440_p1;
wire   [7:0] zext_ln142_213_fu_6444_p1;
wire   [0:0] icmp_ln899_109_fu_6448_p2;
wire   [0:0] xor_ln899_109_fu_6453_p2;
wire  signed [6:0] sext_ln142_41_fu_6463_p1;
wire   [7:0] zext_ln142_215_fu_6467_p1;
wire   [0:0] icmp_ln899_110_fu_6471_p2;
wire   [0:0] xor_ln899_110_fu_6476_p2;
wire  signed [6:0] sext_ln142_42_fu_6486_p1;
wire   [7:0] zext_ln142_217_fu_6490_p1;
wire   [0:0] icmp_ln899_111_fu_6494_p2;
wire   [0:0] xor_ln899_111_fu_6499_p2;
wire  signed [6:0] sext_ln142_43_fu_6509_p1;
wire   [7:0] zext_ln142_219_fu_6513_p1;
wire   [0:0] icmp_ln899_112_fu_6517_p2;
wire   [0:0] xor_ln899_112_fu_6522_p2;
wire  signed [6:0] sext_ln142_44_fu_6532_p1;
wire   [7:0] zext_ln142_221_fu_6536_p1;
wire   [0:0] icmp_ln899_113_fu_6540_p2;
wire   [0:0] xor_ln899_113_fu_6545_p2;
wire  signed [6:0] sext_ln142_45_fu_6555_p1;
wire   [7:0] zext_ln142_223_fu_6559_p1;
wire   [0:0] icmp_ln899_114_fu_6563_p2;
wire   [0:0] xor_ln899_114_fu_6568_p2;
wire  signed [6:0] sext_ln142_46_fu_6578_p1;
wire   [7:0] zext_ln142_225_fu_6582_p1;
wire   [0:0] icmp_ln899_115_fu_6586_p2;
wire   [0:0] xor_ln899_115_fu_6591_p2;
wire  signed [6:0] sext_ln142_47_fu_6601_p1;
wire   [7:0] zext_ln142_227_fu_6605_p1;
wire   [0:0] icmp_ln899_116_fu_6609_p2;
wire   [0:0] xor_ln899_116_fu_6614_p2;
wire  signed [6:0] sext_ln142_48_fu_6624_p1;
wire   [7:0] zext_ln142_229_fu_6628_p1;
wire   [0:0] icmp_ln899_117_fu_6632_p2;
wire   [0:0] xor_ln899_117_fu_6637_p2;
wire  signed [6:0] sext_ln142_49_fu_6647_p1;
wire   [7:0] zext_ln142_231_fu_6651_p1;
wire   [0:0] icmp_ln899_118_fu_6655_p2;
wire   [0:0] xor_ln899_118_fu_6660_p2;
wire  signed [6:0] sext_ln142_50_fu_6670_p1;
wire   [7:0] zext_ln142_233_fu_6674_p1;
wire   [0:0] icmp_ln899_119_fu_6678_p2;
wire   [0:0] xor_ln899_119_fu_6683_p2;
wire  signed [6:0] sext_ln142_51_fu_6693_p1;
wire   [7:0] zext_ln142_235_fu_6697_p1;
wire   [0:0] icmp_ln899_120_fu_6701_p2;
wire   [0:0] xor_ln899_120_fu_6706_p2;
wire  signed [6:0] sext_ln142_52_fu_6716_p1;
wire   [7:0] zext_ln142_237_fu_6720_p1;
wire   [0:0] icmp_ln899_121_fu_6724_p2;
wire   [0:0] xor_ln899_121_fu_6729_p2;
wire  signed [6:0] sext_ln142_53_fu_6739_p1;
wire   [7:0] zext_ln142_239_fu_6743_p1;
wire   [0:0] icmp_ln899_122_fu_6747_p2;
wire   [0:0] xor_ln899_122_fu_6752_p2;
wire  signed [6:0] sext_ln142_54_fu_6762_p1;
wire   [7:0] zext_ln142_241_fu_6766_p1;
wire   [0:0] icmp_ln899_123_fu_6770_p2;
wire   [0:0] xor_ln899_123_fu_6775_p2;
wire  signed [6:0] sext_ln142_55_fu_6785_p1;
wire   [7:0] zext_ln142_243_fu_6789_p1;
wire   [0:0] icmp_ln899_124_fu_6793_p2;
wire   [0:0] xor_ln899_124_fu_6798_p2;
wire  signed [6:0] sext_ln142_56_fu_6808_p1;
wire   [7:0] zext_ln142_245_fu_6812_p1;
wire   [0:0] icmp_ln899_125_fu_6816_p2;
wire   [0:0] xor_ln899_125_fu_6821_p2;
wire   [7:0] select_ln142_5_fu_6831_p3;
wire   [0:0] icmp_ln899_126_fu_6839_p2;
wire   [0:0] xor_ln899_126_fu_6844_p2;
wire   [0:0] icmp_ln899_127_fu_6854_p2;
wire   [0:0] xor_ln899_127_fu_6859_p2;
wire   [0:0] icmp_ln899_128_fu_6869_p2;
wire   [0:0] xor_ln899_128_fu_6874_p2;
wire   [0:0] icmp_ln899_129_fu_6884_p2;
wire   [0:0] xor_ln899_129_fu_6889_p2;
wire   [0:0] icmp_ln899_130_fu_6899_p2;
wire   [0:0] xor_ln899_130_fu_6904_p2;
wire   [0:0] icmp_ln899_131_fu_6914_p2;
wire   [0:0] xor_ln899_131_fu_6919_p2;
wire   [0:0] icmp_ln899_132_fu_6929_p2;
wire   [0:0] xor_ln899_132_fu_6934_p2;
wire   [0:0] icmp_ln899_133_fu_6944_p2;
wire   [0:0] xor_ln899_133_fu_6949_p2;
wire   [0:0] icmp_ln899_134_fu_6959_p2;
wire   [0:0] xor_ln899_134_fu_6964_p2;
wire   [0:0] icmp_ln899_135_fu_6974_p2;
wire   [0:0] xor_ln899_135_fu_6979_p2;
wire   [0:0] icmp_ln899_136_fu_6989_p2;
wire   [0:0] xor_ln899_136_fu_6994_p2;
wire   [0:0] icmp_ln899_137_fu_7004_p2;
wire   [0:0] xor_ln899_137_fu_7009_p2;
wire   [0:0] icmp_ln899_138_fu_7019_p2;
wire   [0:0] xor_ln899_138_fu_7024_p2;
wire   [0:0] icmp_ln899_139_fu_7034_p2;
wire   [0:0] xor_ln899_139_fu_7039_p2;
wire   [0:0] icmp_ln899_140_fu_7049_p2;
wire   [0:0] xor_ln899_140_fu_7054_p2;
wire   [0:0] icmp_ln899_141_fu_7064_p2;
wire   [0:0] xor_ln899_141_fu_7069_p2;
wire   [0:0] icmp_ln899_142_fu_7079_p2;
wire   [0:0] xor_ln899_142_fu_7084_p2;
wire   [0:0] icmp_ln899_143_fu_7094_p2;
wire   [0:0] xor_ln899_143_fu_7099_p2;
wire   [0:0] icmp_ln899_144_fu_7109_p2;
wire   [0:0] xor_ln899_144_fu_7114_p2;
wire   [0:0] icmp_ln899_145_fu_7124_p2;
wire   [0:0] xor_ln899_145_fu_7129_p2;
wire   [0:0] icmp_ln899_146_fu_7139_p2;
wire   [0:0] xor_ln899_146_fu_7144_p2;
wire   [0:0] icmp_ln899_147_fu_7154_p2;
wire   [0:0] xor_ln899_147_fu_7159_p2;
wire   [0:0] icmp_ln899_148_fu_7169_p2;
wire   [0:0] xor_ln899_148_fu_7174_p2;
wire   [0:0] icmp_ln899_149_fu_7184_p2;
wire   [0:0] xor_ln899_149_fu_7189_p2;
wire   [0:0] icmp_ln899_150_fu_7199_p2;
wire   [0:0] xor_ln899_150_fu_7204_p2;
wire   [0:0] icmp_ln899_151_fu_7214_p2;
wire   [0:0] xor_ln899_151_fu_7219_p2;
wire   [0:0] icmp_ln899_152_fu_7229_p2;
wire   [0:0] xor_ln899_152_fu_7234_p2;
wire   [0:0] icmp_ln899_153_fu_7244_p2;
wire   [0:0] xor_ln899_153_fu_7249_p2;
wire   [0:0] icmp_ln899_154_fu_7259_p2;
wire   [0:0] xor_ln899_154_fu_7264_p2;
wire   [0:0] icmp_ln899_155_fu_7274_p2;
wire   [0:0] xor_ln899_155_fu_7279_p2;
wire   [0:0] icmp_ln899_156_fu_7289_p2;
wire   [0:0] xor_ln899_156_fu_7294_p2;
wire   [0:0] icmp_ln899_157_fu_7304_p2;
wire   [0:0] xor_ln899_157_fu_7309_p2;
wire   [0:0] icmp_ln899_158_fu_7319_p2;
wire   [0:0] xor_ln899_158_fu_7324_p2;
wire   [0:0] icmp_ln899_159_fu_7334_p2;
wire   [0:0] xor_ln899_159_fu_7339_p2;
wire   [0:0] icmp_ln899_160_fu_7349_p2;
wire   [0:0] xor_ln899_160_fu_7354_p2;
wire   [0:0] icmp_ln899_161_fu_7364_p2;
wire   [0:0] xor_ln899_161_fu_7369_p2;
wire   [0:0] icmp_ln899_162_fu_7379_p2;
wire   [0:0] xor_ln899_162_fu_7384_p2;
wire   [0:0] icmp_ln899_163_fu_7394_p2;
wire   [0:0] xor_ln899_163_fu_7399_p2;
wire   [0:0] icmp_ln899_164_fu_7409_p2;
wire   [0:0] xor_ln899_164_fu_7414_p2;
wire   [0:0] icmp_ln899_165_fu_7424_p2;
wire   [0:0] xor_ln899_165_fu_7429_p2;
wire   [0:0] icmp_ln899_166_fu_7439_p2;
wire   [0:0] xor_ln899_166_fu_7444_p2;
wire   [0:0] icmp_ln899_167_fu_7454_p2;
wire   [0:0] xor_ln899_167_fu_7459_p2;
wire   [0:0] icmp_ln899_168_fu_7469_p2;
wire   [0:0] xor_ln899_168_fu_7474_p2;
wire   [0:0] icmp_ln899_169_fu_7484_p2;
wire   [0:0] xor_ln899_169_fu_7489_p2;
wire   [0:0] icmp_ln899_170_fu_7499_p2;
wire   [0:0] xor_ln899_170_fu_7504_p2;
wire   [0:0] icmp_ln899_171_fu_7514_p2;
wire   [0:0] xor_ln899_171_fu_7519_p2;
wire   [0:0] icmp_ln899_172_fu_7529_p2;
wire   [0:0] xor_ln899_172_fu_7534_p2;
wire   [0:0] icmp_ln899_173_fu_7544_p2;
wire   [0:0] xor_ln899_173_fu_7549_p2;
wire   [0:0] icmp_ln899_174_fu_7559_p2;
wire   [0:0] xor_ln899_174_fu_7564_p2;
wire   [0:0] icmp_ln899_175_fu_7574_p2;
wire   [0:0] xor_ln899_175_fu_7579_p2;
wire   [0:0] icmp_ln899_176_fu_7589_p2;
wire   [0:0] xor_ln899_176_fu_7594_p2;
wire   [0:0] icmp_ln899_177_fu_7604_p2;
wire   [0:0] xor_ln899_177_fu_7609_p2;
wire   [0:0] icmp_ln899_178_fu_7619_p2;
wire   [0:0] xor_ln899_178_fu_7624_p2;
wire   [0:0] icmp_ln899_179_fu_7634_p2;
wire   [0:0] xor_ln899_179_fu_7639_p2;
wire   [0:0] icmp_ln899_180_fu_7649_p2;
wire   [0:0] xor_ln899_180_fu_7654_p2;
wire   [0:0] icmp_ln899_181_fu_7664_p2;
wire   [0:0] xor_ln899_181_fu_7669_p2;
wire   [0:0] icmp_ln899_182_fu_7679_p2;
wire   [0:0] xor_ln899_182_fu_7684_p2;
wire   [0:0] icmp_ln899_183_fu_7694_p2;
wire   [0:0] xor_ln899_183_fu_7699_p2;
wire   [0:0] icmp_ln899_184_fu_7709_p2;
wire   [0:0] xor_ln899_184_fu_7714_p2;
wire   [0:0] icmp_ln899_185_fu_7724_p2;
wire   [0:0] xor_ln899_185_fu_7729_p2;
wire   [0:0] icmp_ln899_186_fu_7739_p2;
wire   [0:0] xor_ln899_186_fu_7744_p2;
wire   [0:0] icmp_ln899_187_fu_7754_p2;
wire   [0:0] xor_ln899_187_fu_7759_p2;
wire   [0:0] icmp_ln899_188_fu_7769_p2;
wire   [0:0] xor_ln899_188_fu_7774_p2;
wire   [0:0] icmp_ln899_189_fu_7784_p2;
wire   [0:0] xor_ln899_189_fu_7789_p2;
wire   [0:0] icmp_ln899_190_fu_7799_p2;
wire   [0:0] xor_ln899_190_fu_7804_p2;
wire   [0:0] icmp_ln899_191_fu_7814_p2;
wire   [0:0] xor_ln899_191_fu_7819_p2;
wire  signed [7:0] sext_ln142_57_fu_7829_p1;
wire   [0:0] icmp_ln899_192_fu_7833_p2;
wire   [0:0] xor_ln899_192_fu_7838_p2;
wire  signed [7:0] sext_ln142_58_fu_7848_p1;
wire   [0:0] icmp_ln899_193_fu_7852_p2;
wire   [0:0] xor_ln899_193_fu_7857_p2;
wire  signed [7:0] sext_ln142_59_fu_7867_p1;
wire   [0:0] icmp_ln899_194_fu_7871_p2;
wire   [0:0] xor_ln899_194_fu_7876_p2;
wire  signed [7:0] sext_ln142_60_fu_7886_p1;
wire   [0:0] icmp_ln899_195_fu_7890_p2;
wire   [0:0] xor_ln899_195_fu_7895_p2;
wire  signed [7:0] sext_ln142_61_fu_7905_p1;
wire   [0:0] icmp_ln899_196_fu_7909_p2;
wire   [0:0] xor_ln899_196_fu_7914_p2;
wire  signed [7:0] sext_ln142_62_fu_7924_p1;
wire   [0:0] icmp_ln899_197_fu_7928_p2;
wire   [0:0] xor_ln899_197_fu_7933_p2;
wire  signed [7:0] sext_ln142_63_fu_7943_p1;
wire   [0:0] icmp_ln899_198_fu_7947_p2;
wire   [0:0] xor_ln899_198_fu_7952_p2;
wire  signed [7:0] sext_ln142_64_fu_7962_p1;
wire   [0:0] icmp_ln899_199_fu_7966_p2;
wire   [0:0] xor_ln899_199_fu_7971_p2;
wire  signed [7:0] sext_ln142_65_fu_7981_p1;
wire   [0:0] icmp_ln899_200_fu_7985_p2;
wire   [0:0] xor_ln899_200_fu_7990_p2;
wire  signed [7:0] sext_ln142_66_fu_8000_p1;
wire   [0:0] icmp_ln899_201_fu_8004_p2;
wire   [0:0] xor_ln899_201_fu_8009_p2;
wire  signed [7:0] sext_ln142_67_fu_8019_p1;
wire   [0:0] icmp_ln899_202_fu_8023_p2;
wire   [0:0] xor_ln899_202_fu_8028_p2;
wire  signed [7:0] sext_ln142_68_fu_8038_p1;
wire   [0:0] icmp_ln899_203_fu_8042_p2;
wire   [0:0] xor_ln899_203_fu_8047_p2;
wire  signed [7:0] sext_ln142_69_fu_8057_p1;
wire   [0:0] icmp_ln899_204_fu_8061_p2;
wire   [0:0] xor_ln899_204_fu_8066_p2;
wire  signed [7:0] sext_ln142_70_fu_8076_p1;
wire   [0:0] icmp_ln899_205_fu_8080_p2;
wire   [0:0] xor_ln899_205_fu_8085_p2;
wire  signed [7:0] sext_ln142_71_fu_8095_p1;
wire   [0:0] icmp_ln899_206_fu_8099_p2;
wire   [0:0] xor_ln899_206_fu_8104_p2;
wire  signed [7:0] sext_ln142_72_fu_8114_p1;
wire   [0:0] icmp_ln899_207_fu_8118_p2;
wire   [0:0] xor_ln899_207_fu_8123_p2;
wire  signed [7:0] sext_ln142_73_fu_8133_p1;
wire   [0:0] icmp_ln899_208_fu_8137_p2;
wire   [0:0] xor_ln899_208_fu_8142_p2;
wire  signed [7:0] sext_ln142_74_fu_8152_p1;
wire   [0:0] icmp_ln899_209_fu_8156_p2;
wire   [0:0] xor_ln899_209_fu_8161_p2;
wire  signed [7:0] sext_ln142_75_fu_8171_p1;
wire   [0:0] icmp_ln899_210_fu_8175_p2;
wire   [0:0] xor_ln899_210_fu_8180_p2;
wire  signed [7:0] sext_ln142_76_fu_8190_p1;
wire   [0:0] icmp_ln899_211_fu_8194_p2;
wire   [0:0] xor_ln899_211_fu_8199_p2;
wire  signed [7:0] sext_ln142_77_fu_8209_p1;
wire   [0:0] icmp_ln899_212_fu_8213_p2;
wire   [0:0] xor_ln899_212_fu_8218_p2;
wire  signed [7:0] sext_ln142_78_fu_8228_p1;
wire   [0:0] icmp_ln899_213_fu_8232_p2;
wire   [0:0] xor_ln899_213_fu_8237_p2;
wire  signed [7:0] sext_ln142_79_fu_8247_p1;
wire   [0:0] icmp_ln899_214_fu_8251_p2;
wire   [0:0] xor_ln899_214_fu_8256_p2;
wire  signed [7:0] sext_ln142_80_fu_8266_p1;
wire   [0:0] icmp_ln899_215_fu_8270_p2;
wire   [0:0] xor_ln899_215_fu_8275_p2;
wire  signed [7:0] sext_ln142_81_fu_8285_p1;
wire   [0:0] icmp_ln899_216_fu_8289_p2;
wire   [0:0] xor_ln899_216_fu_8294_p2;
wire  signed [7:0] sext_ln142_82_fu_8304_p1;
wire   [0:0] icmp_ln899_217_fu_8308_p2;
wire   [0:0] xor_ln899_217_fu_8313_p2;
wire  signed [7:0] sext_ln142_83_fu_8323_p1;
wire   [0:0] icmp_ln899_218_fu_8327_p2;
wire   [0:0] xor_ln899_218_fu_8332_p2;
wire  signed [7:0] sext_ln142_84_fu_8342_p1;
wire   [0:0] icmp_ln899_219_fu_8346_p2;
wire   [0:0] xor_ln899_219_fu_8351_p2;
wire  signed [7:0] sext_ln142_85_fu_8361_p1;
wire   [0:0] icmp_ln899_220_fu_8365_p2;
wire   [0:0] xor_ln899_220_fu_8370_p2;
wire  signed [7:0] sext_ln142_86_fu_8380_p1;
wire   [0:0] icmp_ln899_221_fu_8384_p2;
wire   [0:0] xor_ln899_221_fu_8389_p2;
wire  signed [7:0] sext_ln142_87_fu_8399_p1;
wire   [0:0] icmp_ln899_222_fu_8403_p2;
wire   [0:0] xor_ln899_222_fu_8408_p2;
wire  signed [7:0] sext_ln142_88_fu_8418_p1;
wire   [0:0] icmp_ln899_223_fu_8422_p2;
wire   [0:0] xor_ln899_223_fu_8427_p2;
wire  signed [7:0] sext_ln142_89_fu_8437_p1;
wire   [0:0] icmp_ln899_224_fu_8441_p2;
wire   [0:0] xor_ln899_224_fu_8446_p2;
wire  signed [7:0] sext_ln142_90_fu_8456_p1;
wire   [0:0] icmp_ln899_225_fu_8460_p2;
wire   [0:0] xor_ln899_225_fu_8465_p2;
wire  signed [7:0] sext_ln142_91_fu_8475_p1;
wire   [0:0] icmp_ln899_226_fu_8479_p2;
wire   [0:0] xor_ln899_226_fu_8484_p2;
wire  signed [7:0] sext_ln142_92_fu_8494_p1;
wire   [0:0] icmp_ln899_227_fu_8498_p2;
wire   [0:0] xor_ln899_227_fu_8503_p2;
wire  signed [7:0] sext_ln142_93_fu_8513_p1;
wire   [0:0] icmp_ln899_228_fu_8517_p2;
wire   [0:0] xor_ln899_228_fu_8522_p2;
wire  signed [7:0] sext_ln142_94_fu_8532_p1;
wire   [0:0] icmp_ln899_229_fu_8536_p2;
wire   [0:0] xor_ln899_229_fu_8541_p2;
wire  signed [7:0] sext_ln142_95_fu_8551_p1;
wire   [0:0] icmp_ln899_230_fu_8555_p2;
wire   [0:0] xor_ln899_230_fu_8560_p2;
wire  signed [7:0] sext_ln142_96_fu_8570_p1;
wire   [0:0] icmp_ln899_231_fu_8574_p2;
wire   [0:0] xor_ln899_231_fu_8579_p2;
wire  signed [7:0] sext_ln142_97_fu_8589_p1;
wire   [0:0] icmp_ln899_232_fu_8593_p2;
wire   [0:0] xor_ln899_232_fu_8598_p2;
wire  signed [7:0] sext_ln142_98_fu_8608_p1;
wire   [0:0] icmp_ln899_233_fu_8612_p2;
wire   [0:0] xor_ln899_233_fu_8617_p2;
wire  signed [7:0] sext_ln142_99_fu_8627_p1;
wire   [0:0] icmp_ln899_234_fu_8631_p2;
wire   [0:0] xor_ln899_234_fu_8636_p2;
wire  signed [7:0] sext_ln142_100_fu_8646_p1;
wire   [0:0] icmp_ln899_235_fu_8650_p2;
wire   [0:0] xor_ln899_235_fu_8655_p2;
wire  signed [7:0] sext_ln142_101_fu_8665_p1;
wire   [0:0] icmp_ln899_236_fu_8669_p2;
wire   [0:0] xor_ln899_236_fu_8674_p2;
wire  signed [7:0] sext_ln142_102_fu_8684_p1;
wire   [0:0] icmp_ln899_237_fu_8688_p2;
wire   [0:0] xor_ln899_237_fu_8693_p2;
wire  signed [7:0] sext_ln142_103_fu_8703_p1;
wire   [0:0] icmp_ln899_238_fu_8707_p2;
wire   [0:0] xor_ln899_238_fu_8712_p2;
wire  signed [7:0] sext_ln142_104_fu_8722_p1;
wire   [0:0] icmp_ln899_239_fu_8726_p2;
wire   [0:0] xor_ln899_239_fu_8731_p2;
wire  signed [7:0] sext_ln142_105_fu_8741_p1;
wire   [0:0] icmp_ln899_240_fu_8745_p2;
wire   [0:0] xor_ln899_240_fu_8750_p2;
wire  signed [7:0] sext_ln142_106_fu_8760_p1;
wire   [0:0] icmp_ln899_241_fu_8764_p2;
wire   [0:0] xor_ln899_241_fu_8769_p2;
wire  signed [7:0] sext_ln142_107_fu_8779_p1;
wire   [0:0] icmp_ln899_242_fu_8783_p2;
wire   [0:0] xor_ln899_242_fu_8788_p2;
wire  signed [7:0] sext_ln142_108_fu_8798_p1;
wire   [0:0] icmp_ln899_243_fu_8802_p2;
wire   [0:0] xor_ln899_243_fu_8807_p2;
wire  signed [7:0] sext_ln142_109_fu_8817_p1;
wire   [0:0] icmp_ln899_244_fu_8821_p2;
wire   [0:0] xor_ln899_244_fu_8826_p2;
wire  signed [7:0] sext_ln142_110_fu_8836_p1;
wire   [0:0] icmp_ln899_245_fu_8840_p2;
wire   [0:0] xor_ln899_245_fu_8845_p2;
wire  signed [7:0] sext_ln142_111_fu_8855_p1;
wire   [0:0] icmp_ln899_246_fu_8859_p2;
wire   [0:0] xor_ln899_246_fu_8864_p2;
wire  signed [7:0] sext_ln142_112_fu_8874_p1;
wire   [0:0] icmp_ln899_247_fu_8878_p2;
wire   [0:0] xor_ln899_247_fu_8883_p2;
wire  signed [7:0] sext_ln142_113_fu_8893_p1;
wire   [0:0] icmp_ln899_248_fu_8897_p2;
wire   [0:0] xor_ln899_248_fu_8902_p2;
wire  signed [7:0] sext_ln142_114_fu_8912_p1;
wire   [0:0] icmp_ln899_249_fu_8916_p2;
wire   [0:0] xor_ln899_249_fu_8921_p2;
wire  signed [7:0] sext_ln142_115_fu_8931_p1;
wire   [0:0] icmp_ln899_250_fu_8935_p2;
wire   [0:0] xor_ln899_250_fu_8940_p2;
wire  signed [7:0] sext_ln142_116_fu_8950_p1;
wire   [0:0] icmp_ln899_251_fu_8954_p2;
wire   [0:0] xor_ln899_251_fu_8959_p2;
wire  signed [7:0] sext_ln142_117_fu_8969_p1;
wire   [0:0] icmp_ln899_252_fu_8973_p2;
wire   [0:0] xor_ln899_252_fu_8978_p2;
wire  signed [7:0] sext_ln142_118_fu_8988_p1;
wire   [0:0] icmp_ln899_253_fu_8992_p2;
wire   [0:0] xor_ln899_253_fu_8997_p2;
wire  signed [7:0] sext_ln142_119_fu_9007_p1;
wire   [0:0] icmp_ln899_254_fu_9011_p2;
wire   [0:0] xor_ln899_254_fu_9016_p2;
wire   [1:0] zext_ln142_6_fu_4265_p1;
wire   [1:0] zext_ln142_8_fu_4284_p1;
wire   [1:0] add_ln700_2_fu_9026_p2;
wire   [1:0] zext_ln142_10_fu_4307_p1;
wire   [1:0] zext_ln142_11_fu_4330_p1;
wire   [1:0] add_ln700_3_fu_9036_p2;
wire   [2:0] zext_ln700_3_fu_9042_p1;
wire   [2:0] zext_ln700_2_fu_9032_p1;
wire   [1:0] zext_ln142_13_fu_4349_p1;
wire   [1:0] zext_ln142_15_fu_4368_p1;
wire   [1:0] add_ln700_6_fu_9052_p2;
wire   [1:0] zext_ln142_17_fu_4387_p1;
wire   [1:0] zext_ln142_19_fu_4406_p1;
wire   [1:0] add_ln700_7_fu_9062_p2;
wire   [2:0] zext_ln700_6_fu_9068_p1;
wire   [2:0] zext_ln700_5_fu_9058_p1;
wire   [1:0] zext_ln142_21_fu_4429_p1;
wire   [1:0] zext_ln142_23_fu_4452_p1;
wire   [1:0] add_ln700_9_fu_9078_p2;
wire   [1:0] zext_ln142_25_fu_4475_p1;
wire   [1:0] zext_ln142_26_fu_4498_p1;
wire   [1:0] add_ln700_10_fu_9088_p2;
wire   [2:0] zext_ln700_9_fu_9094_p1;
wire   [2:0] zext_ln700_8_fu_9084_p1;
wire   [1:0] zext_ln142_28_fu_4517_p1;
wire   [1:0] zext_ln142_30_fu_4536_p1;
wire   [1:0] add_ln700_14_fu_9104_p2;
wire   [1:0] zext_ln142_32_fu_4555_p1;
wire   [1:0] zext_ln142_34_fu_4574_p1;
wire   [1:0] add_ln700_15_fu_9114_p2;
wire   [2:0] zext_ln700_13_fu_9120_p1;
wire   [2:0] zext_ln700_12_fu_9110_p1;
wire   [1:0] zext_ln142_36_fu_4593_p1;
wire   [1:0] zext_ln142_38_fu_4612_p1;
wire   [1:0] add_ln700_17_fu_9130_p2;
wire   [1:0] zext_ln142_40_fu_4631_p1;
wire   [1:0] zext_ln142_42_fu_4650_p1;
wire   [1:0] add_ln700_18_fu_9140_p2;
wire   [2:0] zext_ln700_16_fu_9146_p1;
wire   [2:0] zext_ln700_15_fu_9136_p1;
wire   [1:0] zext_ln142_44_fu_4673_p1;
wire   [1:0] zext_ln142_46_fu_4696_p1;
wire   [1:0] add_ln700_21_fu_9156_p2;
wire   [1:0] zext_ln142_48_fu_4719_p1;
wire   [1:0] zext_ln142_50_fu_4742_p1;
wire   [1:0] add_ln700_22_fu_9166_p2;
wire   [2:0] zext_ln700_20_fu_9172_p1;
wire   [2:0] zext_ln700_19_fu_9162_p1;
wire   [1:0] zext_ln142_52_fu_4765_p1;
wire   [1:0] zext_ln142_54_fu_4788_p1;
wire   [1:0] add_ln700_24_fu_9182_p2;
wire   [1:0] zext_ln142_56_fu_4811_p1;
wire   [1:0] zext_ln142_57_fu_4834_p1;
wire   [1:0] add_ln700_25_fu_9192_p2;
wire   [2:0] zext_ln700_23_fu_9198_p1;
wire   [2:0] zext_ln700_22_fu_9188_p1;
wire   [1:0] zext_ln142_59_fu_4853_p1;
wire   [1:0] zext_ln142_61_fu_4872_p1;
wire   [1:0] add_ln700_30_fu_9208_p2;
wire   [1:0] zext_ln142_63_fu_4891_p1;
wire   [1:0] zext_ln142_65_fu_4910_p1;
wire   [1:0] add_ln700_31_fu_9218_p2;
wire   [2:0] zext_ln700_28_fu_9224_p1;
wire   [2:0] zext_ln700_27_fu_9214_p1;
wire   [1:0] zext_ln142_67_fu_4929_p1;
wire   [1:0] zext_ln142_69_fu_4948_p1;
wire   [1:0] add_ln700_33_fu_9234_p2;
wire   [1:0] zext_ln142_71_fu_4967_p1;
wire   [1:0] zext_ln142_73_fu_4986_p1;
wire   [1:0] add_ln700_34_fu_9244_p2;
wire   [2:0] zext_ln700_31_fu_9250_p1;
wire   [2:0] zext_ln700_30_fu_9240_p1;
wire   [1:0] zext_ln142_75_fu_5005_p1;
wire   [1:0] zext_ln142_77_fu_5024_p1;
wire   [1:0] add_ln700_37_fu_9260_p2;
wire   [1:0] zext_ln142_79_fu_5043_p1;
wire   [1:0] zext_ln142_81_fu_5062_p1;
wire   [1:0] add_ln700_38_fu_9270_p2;
wire   [2:0] zext_ln700_35_fu_9276_p1;
wire   [2:0] zext_ln700_34_fu_9266_p1;
wire   [1:0] zext_ln142_83_fu_5081_p1;
wire   [1:0] zext_ln142_85_fu_5100_p1;
wire   [1:0] add_ln700_40_fu_9286_p2;
wire   [1:0] zext_ln142_87_fu_5119_p1;
wire   [1:0] zext_ln142_89_fu_5138_p1;
wire   [1:0] add_ln700_41_fu_9296_p2;
wire   [2:0] zext_ln700_38_fu_9302_p1;
wire   [2:0] zext_ln700_37_fu_9292_p1;
wire   [1:0] zext_ln142_91_fu_5161_p1;
wire   [1:0] zext_ln142_93_fu_5184_p1;
wire   [1:0] add_ln700_45_fu_9312_p2;
wire   [1:0] zext_ln142_95_fu_5207_p1;
wire   [1:0] zext_ln142_97_fu_5230_p1;
wire   [1:0] add_ln700_46_fu_9322_p2;
wire   [2:0] zext_ln700_43_fu_9328_p1;
wire   [2:0] zext_ln700_42_fu_9318_p1;
wire   [1:0] zext_ln142_99_fu_5253_p1;
wire   [1:0] zext_ln142_101_fu_5276_p1;
wire   [1:0] add_ln700_48_fu_9338_p2;
wire   [1:0] zext_ln142_103_fu_5299_p1;
wire   [1:0] zext_ln142_105_fu_5322_p1;
wire   [1:0] add_ln700_49_fu_9348_p2;
wire   [2:0] zext_ln700_46_fu_9354_p1;
wire   [2:0] zext_ln700_45_fu_9344_p1;
wire   [1:0] zext_ln142_107_fu_5345_p1;
wire   [1:0] zext_ln142_109_fu_5368_p1;
wire   [1:0] add_ln700_52_fu_9364_p2;
wire   [1:0] zext_ln142_111_fu_5391_p1;
wire   [1:0] zext_ln142_113_fu_5414_p1;
wire   [1:0] add_ln700_53_fu_9374_p2;
wire   [2:0] zext_ln700_50_fu_9380_p1;
wire   [2:0] zext_ln700_49_fu_9370_p1;
wire   [1:0] zext_ln142_115_fu_5437_p1;
wire   [1:0] zext_ln142_117_fu_5460_p1;
wire   [1:0] add_ln700_55_fu_9390_p2;
wire   [1:0] zext_ln142_119_fu_5483_p1;
wire   [1:0] zext_ln142_120_fu_5506_p1;
wire   [1:0] add_ln700_56_fu_9400_p2;
wire   [2:0] zext_ln700_53_fu_9406_p1;
wire   [2:0] zext_ln700_52_fu_9396_p1;
wire   [1:0] zext_ln142_122_fu_5525_p1;
wire   [1:0] zext_ln142_124_fu_5544_p1;
wire   [1:0] add_ln700_62_fu_9416_p2;
wire   [1:0] zext_ln142_126_fu_5563_p1;
wire   [1:0] zext_ln142_128_fu_5582_p1;
wire   [1:0] add_ln700_63_fu_9426_p2;
wire   [2:0] zext_ln700_59_fu_9432_p1;
wire   [2:0] zext_ln700_58_fu_9422_p1;
wire   [1:0] zext_ln142_130_fu_5601_p1;
wire   [1:0] zext_ln142_132_fu_5620_p1;
wire   [1:0] add_ln700_65_fu_9442_p2;
wire   [1:0] zext_ln142_134_fu_5639_p1;
wire   [1:0] zext_ln142_136_fu_5658_p1;
wire   [1:0] add_ln700_66_fu_9452_p2;
wire   [2:0] zext_ln700_62_fu_9458_p1;
wire   [2:0] zext_ln700_61_fu_9448_p1;
wire   [1:0] zext_ln142_138_fu_5677_p1;
wire   [1:0] zext_ln142_140_fu_5696_p1;
wire   [1:0] add_ln700_69_fu_9468_p2;
wire   [1:0] zext_ln142_142_fu_5715_p1;
wire   [1:0] zext_ln142_144_fu_5734_p1;
wire   [1:0] add_ln700_70_fu_9478_p2;
wire   [2:0] zext_ln700_66_fu_9484_p1;
wire   [2:0] zext_ln700_65_fu_9474_p1;
wire   [1:0] zext_ln142_146_fu_5753_p1;
wire   [1:0] zext_ln142_148_fu_5772_p1;
wire   [1:0] add_ln700_72_fu_9494_p2;
wire   [1:0] zext_ln142_150_fu_5791_p1;
wire   [1:0] zext_ln142_152_fu_5810_p1;
wire   [1:0] add_ln700_73_fu_9504_p2;
wire   [2:0] zext_ln700_69_fu_9510_p1;
wire   [2:0] zext_ln700_68_fu_9500_p1;
wire   [1:0] zext_ln142_154_fu_5829_p1;
wire   [1:0] zext_ln142_156_fu_5848_p1;
wire   [1:0] add_ln700_77_fu_9520_p2;
wire   [1:0] zext_ln142_158_fu_5867_p1;
wire   [1:0] zext_ln142_160_fu_5886_p1;
wire   [1:0] add_ln700_78_fu_9530_p2;
wire   [2:0] zext_ln700_74_fu_9536_p1;
wire   [2:0] zext_ln700_73_fu_9526_p1;
wire   [1:0] zext_ln142_162_fu_5905_p1;
wire   [1:0] zext_ln142_164_fu_5924_p1;
wire   [1:0] add_ln700_80_fu_9546_p2;
wire   [1:0] zext_ln142_166_fu_5943_p1;
wire   [1:0] zext_ln142_168_fu_5962_p1;
wire   [1:0] add_ln700_81_fu_9556_p2;
wire   [2:0] zext_ln700_77_fu_9562_p1;
wire   [2:0] zext_ln700_76_fu_9552_p1;
wire   [1:0] zext_ln142_170_fu_5981_p1;
wire   [1:0] zext_ln142_172_fu_6000_p1;
wire   [1:0] add_ln700_84_fu_9572_p2;
wire   [1:0] zext_ln142_174_fu_6019_p1;
wire   [1:0] zext_ln142_176_fu_6038_p1;
wire   [1:0] add_ln700_85_fu_9582_p2;
wire   [2:0] zext_ln700_81_fu_9588_p1;
wire   [2:0] zext_ln700_80_fu_9578_p1;
wire   [1:0] zext_ln142_178_fu_6057_p1;
wire   [1:0] zext_ln142_180_fu_6076_p1;
wire   [1:0] add_ln700_87_fu_9598_p2;
wire   [1:0] zext_ln142_182_fu_6095_p1;
wire   [1:0] zext_ln142_184_fu_6114_p1;
wire   [1:0] add_ln700_88_fu_9608_p2;
wire   [2:0] zext_ln700_84_fu_9614_p1;
wire   [2:0] zext_ln700_83_fu_9604_p1;
wire   [1:0] zext_ln142_186_fu_6137_p1;
wire   [1:0] zext_ln142_188_fu_6160_p1;
wire   [1:0] add_ln700_93_fu_9624_p2;
wire   [1:0] zext_ln142_190_fu_6183_p1;
wire   [1:0] zext_ln142_192_fu_6206_p1;
wire   [1:0] add_ln700_94_fu_9634_p2;
wire   [2:0] zext_ln700_90_fu_9640_p1;
wire   [2:0] zext_ln700_89_fu_9630_p1;
wire   [1:0] zext_ln142_194_fu_6229_p1;
wire   [1:0] zext_ln142_196_fu_6252_p1;
wire   [1:0] add_ln700_96_fu_9650_p2;
wire   [1:0] zext_ln142_198_fu_6275_p1;
wire   [1:0] zext_ln142_200_fu_6298_p1;
wire   [1:0] add_ln700_97_fu_9660_p2;
wire   [2:0] zext_ln700_93_fu_9666_p1;
wire   [2:0] zext_ln700_92_fu_9656_p1;
wire   [1:0] zext_ln142_202_fu_6321_p1;
wire   [1:0] zext_ln142_204_fu_6344_p1;
wire   [1:0] add_ln700_100_fu_9676_p2;
wire   [1:0] zext_ln142_206_fu_6367_p1;
wire   [1:0] zext_ln142_208_fu_6390_p1;
wire   [1:0] add_ln700_101_fu_9686_p2;
wire   [2:0] zext_ln700_97_fu_9692_p1;
wire   [2:0] zext_ln700_96_fu_9682_p1;
wire   [1:0] zext_ln142_210_fu_6413_p1;
wire   [1:0] zext_ln142_212_fu_6436_p1;
wire   [1:0] add_ln700_103_fu_9702_p2;
wire   [1:0] zext_ln142_214_fu_6459_p1;
wire   [1:0] zext_ln142_216_fu_6482_p1;
wire   [1:0] add_ln700_104_fu_9712_p2;
wire   [2:0] zext_ln700_100_fu_9718_p1;
wire   [2:0] zext_ln700_99_fu_9708_p1;
wire   [1:0] zext_ln142_218_fu_6505_p1;
wire   [1:0] zext_ln142_220_fu_6528_p1;
wire   [1:0] add_ln700_108_fu_9728_p2;
wire   [1:0] zext_ln142_222_fu_6551_p1;
wire   [1:0] zext_ln142_224_fu_6574_p1;
wire   [1:0] add_ln700_109_fu_9738_p2;
wire   [2:0] zext_ln700_105_fu_9744_p1;
wire   [2:0] zext_ln700_104_fu_9734_p1;
wire   [1:0] zext_ln142_226_fu_6597_p1;
wire   [1:0] zext_ln142_228_fu_6620_p1;
wire   [1:0] add_ln700_111_fu_9754_p2;
wire   [1:0] zext_ln142_230_fu_6643_p1;
wire   [1:0] zext_ln142_232_fu_6666_p1;
wire   [1:0] add_ln700_112_fu_9764_p2;
wire   [2:0] zext_ln700_108_fu_9770_p1;
wire   [2:0] zext_ln700_107_fu_9760_p1;
wire   [1:0] zext_ln142_234_fu_6689_p1;
wire   [1:0] zext_ln142_236_fu_6712_p1;
wire   [1:0] add_ln700_115_fu_9780_p2;
wire   [1:0] zext_ln142_238_fu_6735_p1;
wire   [1:0] zext_ln142_240_fu_6758_p1;
wire   [1:0] add_ln700_116_fu_9790_p2;
wire   [2:0] zext_ln700_112_fu_9796_p1;
wire   [2:0] zext_ln700_111_fu_9786_p1;
wire   [1:0] zext_ln142_242_fu_6781_p1;
wire   [1:0] zext_ln142_244_fu_6804_p1;
wire   [1:0] add_ln700_118_fu_9806_p2;
wire   [1:0] zext_ln142_246_fu_6827_p1;
wire   [1:0] zext_ln142_247_fu_6850_p1;
wire   [1:0] add_ln700_119_fu_9816_p2;
wire   [2:0] zext_ln700_115_fu_9822_p1;
wire   [2:0] zext_ln700_114_fu_9812_p1;
wire   [1:0] zext_ln142_248_fu_6865_p1;
wire   [1:0] zext_ln142_249_fu_6880_p1;
wire   [1:0] add_ln700_126_fu_9832_p2;
wire   [1:0] zext_ln142_250_fu_6895_p1;
wire   [1:0] zext_ln142_251_fu_6910_p1;
wire   [1:0] add_ln700_127_fu_9842_p2;
wire   [2:0] zext_ln700_122_fu_9848_p1;
wire   [2:0] zext_ln700_121_fu_9838_p1;
wire   [1:0] zext_ln142_252_fu_6925_p1;
wire   [1:0] zext_ln142_253_fu_6940_p1;
wire   [1:0] add_ln700_129_fu_9858_p2;
wire   [1:0] zext_ln142_254_fu_6955_p1;
wire   [1:0] zext_ln142_255_fu_6970_p1;
wire   [1:0] add_ln700_130_fu_9868_p2;
wire   [2:0] zext_ln700_125_fu_9874_p1;
wire   [2:0] zext_ln700_124_fu_9864_p1;
wire   [1:0] zext_ln142_256_fu_6985_p1;
wire   [1:0] zext_ln142_257_fu_7000_p1;
wire   [1:0] add_ln700_133_fu_9884_p2;
wire   [1:0] zext_ln142_258_fu_7015_p1;
wire   [1:0] zext_ln142_259_fu_7030_p1;
wire   [1:0] add_ln700_134_fu_9894_p2;
wire   [2:0] zext_ln700_129_fu_9900_p1;
wire   [2:0] zext_ln700_128_fu_9890_p1;
wire   [1:0] zext_ln142_260_fu_7045_p1;
wire   [1:0] zext_ln142_261_fu_7060_p1;
wire   [1:0] add_ln700_136_fu_9910_p2;
wire   [1:0] zext_ln142_262_fu_7075_p1;
wire   [1:0] zext_ln142_263_fu_7090_p1;
wire   [1:0] add_ln700_137_fu_9920_p2;
wire   [2:0] zext_ln700_132_fu_9926_p1;
wire   [2:0] zext_ln700_131_fu_9916_p1;
wire   [1:0] zext_ln142_264_fu_7105_p1;
wire   [1:0] zext_ln142_265_fu_7120_p1;
wire   [1:0] add_ln700_141_fu_9936_p2;
wire   [1:0] zext_ln142_266_fu_7135_p1;
wire   [1:0] zext_ln142_267_fu_7150_p1;
wire   [1:0] add_ln700_142_fu_9946_p2;
wire   [2:0] zext_ln700_137_fu_9952_p1;
wire   [2:0] zext_ln700_136_fu_9942_p1;
wire   [1:0] zext_ln142_268_fu_7165_p1;
wire   [1:0] zext_ln142_269_fu_7180_p1;
wire   [1:0] add_ln700_144_fu_9962_p2;
wire   [1:0] zext_ln142_270_fu_7195_p1;
wire   [1:0] zext_ln142_271_fu_7210_p1;
wire   [1:0] add_ln700_145_fu_9972_p2;
wire   [2:0] zext_ln700_140_fu_9978_p1;
wire   [2:0] zext_ln700_139_fu_9968_p1;
wire   [1:0] zext_ln142_272_fu_7225_p1;
wire   [1:0] zext_ln142_273_fu_7240_p1;
wire   [1:0] add_ln700_148_fu_9988_p2;
wire   [1:0] zext_ln142_274_fu_7255_p1;
wire   [1:0] zext_ln142_275_fu_7270_p1;
wire   [1:0] add_ln700_149_fu_9998_p2;
wire   [2:0] zext_ln700_144_fu_10004_p1;
wire   [2:0] zext_ln700_143_fu_9994_p1;
wire   [1:0] zext_ln142_276_fu_7285_p1;
wire   [1:0] zext_ln142_277_fu_7300_p1;
wire   [1:0] add_ln700_151_fu_10014_p2;
wire   [1:0] zext_ln142_278_fu_7315_p1;
wire   [1:0] zext_ln142_279_fu_7330_p1;
wire   [1:0] add_ln700_152_fu_10024_p2;
wire   [2:0] zext_ln700_147_fu_10030_p1;
wire   [2:0] zext_ln700_146_fu_10020_p1;
wire   [1:0] zext_ln142_280_fu_7345_p1;
wire   [1:0] zext_ln142_281_fu_7360_p1;
wire   [1:0] add_ln700_157_fu_10040_p2;
wire   [1:0] zext_ln142_282_fu_7375_p1;
wire   [1:0] zext_ln142_283_fu_7390_p1;
wire   [1:0] add_ln700_158_fu_10050_p2;
wire   [2:0] zext_ln700_153_fu_10056_p1;
wire   [2:0] zext_ln700_152_fu_10046_p1;
wire   [1:0] zext_ln142_284_fu_7405_p1;
wire   [1:0] zext_ln142_285_fu_7420_p1;
wire   [1:0] add_ln700_160_fu_10066_p2;
wire   [1:0] zext_ln142_286_fu_7435_p1;
wire   [1:0] zext_ln142_287_fu_7450_p1;
wire   [1:0] add_ln700_161_fu_10076_p2;
wire   [2:0] zext_ln700_156_fu_10082_p1;
wire   [2:0] zext_ln700_155_fu_10072_p1;
wire   [1:0] zext_ln142_288_fu_7465_p1;
wire   [1:0] zext_ln142_289_fu_7480_p1;
wire   [1:0] add_ln700_164_fu_10092_p2;
wire   [1:0] zext_ln142_290_fu_7495_p1;
wire   [1:0] zext_ln142_291_fu_7510_p1;
wire   [1:0] add_ln700_165_fu_10102_p2;
wire   [2:0] zext_ln700_160_fu_10108_p1;
wire   [2:0] zext_ln700_159_fu_10098_p1;
wire   [1:0] zext_ln142_292_fu_7525_p1;
wire   [1:0] zext_ln142_293_fu_7540_p1;
wire   [1:0] add_ln700_167_fu_10118_p2;
wire   [1:0] zext_ln142_294_fu_7555_p1;
wire   [1:0] zext_ln142_295_fu_7570_p1;
wire   [1:0] add_ln700_168_fu_10128_p2;
wire   [2:0] zext_ln700_163_fu_10134_p1;
wire   [2:0] zext_ln700_162_fu_10124_p1;
wire   [1:0] zext_ln142_296_fu_7585_p1;
wire   [1:0] zext_ln142_297_fu_7600_p1;
wire   [1:0] add_ln700_172_fu_10144_p2;
wire   [1:0] zext_ln142_298_fu_7615_p1;
wire   [1:0] zext_ln142_299_fu_7630_p1;
wire   [1:0] add_ln700_173_fu_10154_p2;
wire   [2:0] zext_ln700_168_fu_10160_p1;
wire   [2:0] zext_ln700_167_fu_10150_p1;
wire   [1:0] zext_ln142_300_fu_7645_p1;
wire   [1:0] zext_ln142_301_fu_7660_p1;
wire   [1:0] add_ln700_175_fu_10170_p2;
wire   [1:0] zext_ln142_302_fu_7675_p1;
wire   [1:0] zext_ln142_303_fu_7690_p1;
wire   [1:0] add_ln700_176_fu_10180_p2;
wire   [2:0] zext_ln700_171_fu_10186_p1;
wire   [2:0] zext_ln700_170_fu_10176_p1;
wire   [1:0] zext_ln142_304_fu_7705_p1;
wire   [1:0] zext_ln142_305_fu_7720_p1;
wire   [1:0] add_ln700_179_fu_10196_p2;
wire   [1:0] zext_ln142_306_fu_7735_p1;
wire   [1:0] zext_ln142_307_fu_7750_p1;
wire   [1:0] add_ln700_180_fu_10206_p2;
wire   [2:0] zext_ln700_175_fu_10212_p1;
wire   [2:0] zext_ln700_174_fu_10202_p1;
wire   [1:0] zext_ln142_308_fu_7765_p1;
wire   [1:0] zext_ln142_309_fu_7780_p1;
wire   [1:0] add_ln700_182_fu_10222_p2;
wire   [1:0] zext_ln142_310_fu_7795_p1;
wire   [1:0] zext_ln142_311_fu_7810_p1;
wire   [1:0] add_ln700_183_fu_10232_p2;
wire   [2:0] zext_ln700_178_fu_10238_p1;
wire   [2:0] zext_ln700_177_fu_10228_p1;
wire   [1:0] zext_ln142_312_fu_7825_p1;
wire   [1:0] zext_ln142_313_fu_7844_p1;
wire   [1:0] add_ln700_189_fu_10248_p2;
wire   [1:0] zext_ln142_314_fu_7863_p1;
wire   [1:0] zext_ln142_315_fu_7882_p1;
wire   [1:0] add_ln700_190_fu_10258_p2;
wire   [2:0] zext_ln700_185_fu_10264_p1;
wire   [2:0] zext_ln700_184_fu_10254_p1;
wire   [1:0] zext_ln142_316_fu_7901_p1;
wire   [1:0] zext_ln142_317_fu_7920_p1;
wire   [1:0] add_ln700_192_fu_10274_p2;
wire   [1:0] zext_ln142_318_fu_7939_p1;
wire   [1:0] zext_ln142_319_fu_7958_p1;
wire   [1:0] add_ln700_193_fu_10284_p2;
wire   [2:0] zext_ln700_188_fu_10290_p1;
wire   [2:0] zext_ln700_187_fu_10280_p1;
wire   [1:0] zext_ln142_320_fu_7977_p1;
wire   [1:0] zext_ln142_321_fu_7996_p1;
wire   [1:0] add_ln700_196_fu_10300_p2;
wire   [1:0] zext_ln142_322_fu_8015_p1;
wire   [1:0] zext_ln142_323_fu_8034_p1;
wire   [1:0] add_ln700_197_fu_10310_p2;
wire   [2:0] zext_ln700_192_fu_10316_p1;
wire   [2:0] zext_ln700_191_fu_10306_p1;
wire   [1:0] zext_ln142_324_fu_8053_p1;
wire   [1:0] zext_ln142_325_fu_8072_p1;
wire   [1:0] add_ln700_199_fu_10326_p2;
wire   [1:0] zext_ln142_326_fu_8091_p1;
wire   [1:0] zext_ln142_327_fu_8110_p1;
wire   [1:0] add_ln700_200_fu_10336_p2;
wire   [2:0] zext_ln700_195_fu_10342_p1;
wire   [2:0] zext_ln700_194_fu_10332_p1;
wire   [1:0] zext_ln142_328_fu_8129_p1;
wire   [1:0] zext_ln142_329_fu_8148_p1;
wire   [1:0] add_ln700_204_fu_10352_p2;
wire   [1:0] zext_ln142_330_fu_8167_p1;
wire   [1:0] zext_ln142_331_fu_8186_p1;
wire   [1:0] add_ln700_205_fu_10362_p2;
wire   [2:0] zext_ln700_200_fu_10368_p1;
wire   [2:0] zext_ln700_199_fu_10358_p1;
wire   [1:0] zext_ln142_332_fu_8205_p1;
wire   [1:0] zext_ln142_333_fu_8224_p1;
wire   [1:0] add_ln700_207_fu_10378_p2;
wire   [1:0] zext_ln142_334_fu_8243_p1;
wire   [1:0] zext_ln142_335_fu_8262_p1;
wire   [1:0] add_ln700_208_fu_10388_p2;
wire   [2:0] zext_ln700_203_fu_10394_p1;
wire   [2:0] zext_ln700_202_fu_10384_p1;
wire   [1:0] zext_ln142_336_fu_8281_p1;
wire   [1:0] zext_ln142_337_fu_8300_p1;
wire   [1:0] add_ln700_211_fu_10404_p2;
wire   [1:0] zext_ln142_338_fu_8319_p1;
wire   [1:0] zext_ln142_339_fu_8338_p1;
wire   [1:0] add_ln700_212_fu_10414_p2;
wire   [2:0] zext_ln700_207_fu_10420_p1;
wire   [2:0] zext_ln700_206_fu_10410_p1;
wire   [1:0] zext_ln142_340_fu_8357_p1;
wire   [1:0] zext_ln142_341_fu_8376_p1;
wire   [1:0] add_ln700_214_fu_10430_p2;
wire   [1:0] zext_ln142_342_fu_8395_p1;
wire   [1:0] zext_ln142_343_fu_8414_p1;
wire   [1:0] add_ln700_215_fu_10440_p2;
wire   [2:0] zext_ln700_210_fu_10446_p1;
wire   [2:0] zext_ln700_209_fu_10436_p1;
wire   [1:0] zext_ln142_344_fu_8433_p1;
wire   [1:0] zext_ln142_345_fu_8452_p1;
wire   [1:0] add_ln700_220_fu_10456_p2;
wire   [1:0] zext_ln142_346_fu_8471_p1;
wire   [1:0] zext_ln142_347_fu_8490_p1;
wire   [1:0] add_ln700_221_fu_10466_p2;
wire   [2:0] zext_ln700_216_fu_10472_p1;
wire   [2:0] zext_ln700_215_fu_10462_p1;
wire   [1:0] zext_ln142_348_fu_8509_p1;
wire   [1:0] zext_ln142_349_fu_8528_p1;
wire   [1:0] add_ln700_223_fu_10482_p2;
wire   [1:0] zext_ln142_350_fu_8547_p1;
wire   [1:0] zext_ln142_351_fu_8566_p1;
wire   [1:0] add_ln700_224_fu_10492_p2;
wire   [2:0] zext_ln700_219_fu_10498_p1;
wire   [2:0] zext_ln700_218_fu_10488_p1;
wire   [1:0] zext_ln142_352_fu_8585_p1;
wire   [1:0] zext_ln142_353_fu_8604_p1;
wire   [1:0] add_ln700_227_fu_10508_p2;
wire   [1:0] zext_ln142_354_fu_8623_p1;
wire   [1:0] zext_ln142_355_fu_8642_p1;
wire   [1:0] add_ln700_228_fu_10518_p2;
wire   [2:0] zext_ln700_223_fu_10524_p1;
wire   [2:0] zext_ln700_222_fu_10514_p1;
wire   [1:0] zext_ln142_356_fu_8661_p1;
wire   [1:0] zext_ln142_357_fu_8680_p1;
wire   [1:0] add_ln700_230_fu_10534_p2;
wire   [1:0] zext_ln142_358_fu_8699_p1;
wire   [1:0] zext_ln142_359_fu_8718_p1;
wire   [1:0] add_ln700_231_fu_10544_p2;
wire   [2:0] zext_ln700_226_fu_10550_p1;
wire   [2:0] zext_ln700_225_fu_10540_p1;
wire   [1:0] zext_ln142_360_fu_8737_p1;
wire   [1:0] zext_ln142_361_fu_8756_p1;
wire   [1:0] add_ln700_235_fu_10560_p2;
wire   [1:0] zext_ln142_362_fu_8775_p1;
wire   [1:0] zext_ln142_363_fu_8794_p1;
wire   [1:0] add_ln700_236_fu_10570_p2;
wire   [2:0] zext_ln700_231_fu_10576_p1;
wire   [2:0] zext_ln700_230_fu_10566_p1;
wire   [1:0] zext_ln142_364_fu_8813_p1;
wire   [1:0] zext_ln142_365_fu_8832_p1;
wire   [1:0] add_ln700_238_fu_10586_p2;
wire   [1:0] zext_ln142_366_fu_8851_p1;
wire   [1:0] zext_ln142_367_fu_8870_p1;
wire   [1:0] add_ln700_239_fu_10596_p2;
wire   [2:0] zext_ln700_234_fu_10602_p1;
wire   [2:0] zext_ln700_233_fu_10592_p1;
wire   [1:0] zext_ln142_368_fu_8889_p1;
wire   [1:0] zext_ln142_369_fu_8908_p1;
wire   [1:0] add_ln700_242_fu_10612_p2;
wire   [1:0] zext_ln142_370_fu_8927_p1;
wire   [1:0] zext_ln142_371_fu_8946_p1;
wire   [1:0] add_ln700_243_fu_10622_p2;
wire   [2:0] zext_ln700_238_fu_10628_p1;
wire   [2:0] zext_ln700_237_fu_10618_p1;
wire   [1:0] zext_ln142_372_fu_8965_p1;
wire   [1:0] zext_ln142_373_fu_8984_p1;
wire   [1:0] add_ln700_245_fu_10638_p2;
wire   [1:0] zext_ln142_374_fu_9003_p1;
wire   [1:0] zext_ln700_fu_9022_p1;
wire   [1:0] add_ln700_246_fu_10648_p2;
wire   [2:0] zext_ln700_241_fu_10654_p1;
wire   [2:0] zext_ln700_240_fu_10644_p1;
wire   [0:0] xor_ln899_fu_10664_p2;
wire   [0:0] xor_ln899_1_fu_10677_p2;
wire   [0:0] xor_ln899_2_fu_10686_p2;
wire   [1:0] zext_ln142_3_fu_10682_p1;
wire   [1:0] zext_ln142_4_fu_10691_p1;
wire   [1:0] add_ln700_fu_10695_p2;
wire   [7:0] zext_ln700_1_fu_10701_p1;
wire   [7:0] or_ln_fu_10669_p3;
wire   [7:0] zext_ln700_4_fu_10711_p1;
wire   [7:0] add_ln700_1_fu_10705_p2;
wire   [3:0] zext_ln700_10_fu_10723_p1;
wire   [3:0] zext_ln700_7_fu_10720_p1;
wire   [3:0] add_ln700_12_fu_10726_p2;
wire   [7:0] zext_ln700_11_fu_10732_p1;
wire   [7:0] add_ln700_5_fu_10714_p2;
wire   [3:0] zext_ln700_17_fu_10745_p1;
wire   [3:0] zext_ln700_14_fu_10742_p1;
wire   [3:0] add_ln700_20_fu_10748_p2;
wire   [3:0] zext_ln700_24_fu_10761_p1;
wire   [3:0] zext_ln700_21_fu_10758_p1;
wire   [3:0] add_ln700_27_fu_10764_p2;
wire   [4:0] zext_ln700_25_fu_10770_p1;
wire   [4:0] zext_ln700_18_fu_10754_p1;
wire   [3:0] zext_ln700_32_fu_10783_p1;
wire   [3:0] zext_ln700_29_fu_10780_p1;
wire   [3:0] add_ln700_36_fu_10786_p2;
wire   [3:0] zext_ln700_39_fu_10799_p1;
wire   [3:0] zext_ln700_36_fu_10796_p1;
wire   [3:0] add_ln700_43_fu_10802_p2;
wire   [4:0] zext_ln700_40_fu_10808_p1;
wire   [4:0] zext_ln700_33_fu_10792_p1;
wire   [4:0] add_ln700_44_fu_10812_p2;
wire   [3:0] zext_ln700_47_fu_10825_p1;
wire   [3:0] zext_ln700_44_fu_10822_p1;
wire   [3:0] add_ln700_51_fu_10828_p2;
wire   [3:0] zext_ln700_54_fu_10841_p1;
wire   [3:0] zext_ln700_51_fu_10838_p1;
wire   [3:0] add_ln700_58_fu_10844_p2;
wire   [4:0] zext_ln700_55_fu_10850_p1;
wire   [4:0] zext_ln700_48_fu_10834_p1;
wire   [4:0] add_ln700_59_fu_10854_p2;
wire   [5:0] zext_ln700_56_fu_10860_p1;
wire   [5:0] zext_ln700_41_fu_10818_p1;
wire   [3:0] zext_ln700_63_fu_10873_p1;
wire   [3:0] zext_ln700_60_fu_10870_p1;
wire   [3:0] add_ln700_68_fu_10876_p2;
wire   [3:0] zext_ln700_70_fu_10889_p1;
wire   [3:0] zext_ln700_67_fu_10886_p1;
wire   [3:0] add_ln700_75_fu_10892_p2;
wire   [4:0] zext_ln700_71_fu_10898_p1;
wire   [4:0] zext_ln700_64_fu_10882_p1;
wire   [4:0] add_ln700_76_fu_10902_p2;
wire   [3:0] zext_ln700_78_fu_10915_p1;
wire   [3:0] zext_ln700_75_fu_10912_p1;
wire   [3:0] add_ln700_83_fu_10918_p2;
wire   [3:0] zext_ln700_85_fu_10931_p1;
wire   [3:0] zext_ln700_82_fu_10928_p1;
wire   [3:0] add_ln700_90_fu_10934_p2;
wire   [4:0] zext_ln700_86_fu_10940_p1;
wire   [4:0] zext_ln700_79_fu_10924_p1;
wire   [4:0] add_ln700_91_fu_10944_p2;
wire   [5:0] zext_ln700_87_fu_10950_p1;
wire   [5:0] zext_ln700_72_fu_10908_p1;
wire   [5:0] add_ln700_92_fu_10954_p2;
wire   [3:0] zext_ln700_94_fu_10967_p1;
wire   [3:0] zext_ln700_91_fu_10964_p1;
wire   [3:0] add_ln700_99_fu_10970_p2;
wire   [3:0] zext_ln700_101_fu_10983_p1;
wire   [3:0] zext_ln700_98_fu_10980_p1;
wire   [3:0] add_ln700_106_fu_10986_p2;
wire   [4:0] zext_ln700_102_fu_10992_p1;
wire   [4:0] zext_ln700_95_fu_10976_p1;
wire   [4:0] add_ln700_107_fu_10996_p2;
wire   [3:0] zext_ln700_109_fu_11009_p1;
wire   [3:0] zext_ln700_106_fu_11006_p1;
wire   [3:0] add_ln700_114_fu_11012_p2;
wire   [3:0] zext_ln700_116_fu_11025_p1;
wire   [3:0] zext_ln700_113_fu_11022_p1;
wire   [3:0] add_ln700_121_fu_11028_p2;
wire   [4:0] zext_ln700_117_fu_11034_p1;
wire   [4:0] zext_ln700_110_fu_11018_p1;
wire   [4:0] add_ln700_122_fu_11038_p2;
wire   [5:0] zext_ln700_118_fu_11044_p1;
wire   [5:0] zext_ln700_103_fu_11002_p1;
wire   [5:0] add_ln700_123_fu_11048_p2;
wire   [6:0] zext_ln700_119_fu_11054_p1;
wire   [6:0] zext_ln700_88_fu_10960_p1;
wire   [3:0] zext_ln700_126_fu_11067_p1;
wire   [3:0] zext_ln700_123_fu_11064_p1;
wire   [3:0] add_ln700_132_fu_11070_p2;
wire   [3:0] zext_ln700_133_fu_11083_p1;
wire   [3:0] zext_ln700_130_fu_11080_p1;
wire   [3:0] add_ln700_139_fu_11086_p2;
wire   [4:0] zext_ln700_134_fu_11092_p1;
wire   [4:0] zext_ln700_127_fu_11076_p1;
wire   [4:0] add_ln700_140_fu_11096_p2;
wire   [3:0] zext_ln700_141_fu_11109_p1;
wire   [3:0] zext_ln700_138_fu_11106_p1;
wire   [3:0] add_ln700_147_fu_11112_p2;
wire   [3:0] zext_ln700_148_fu_11125_p1;
wire   [3:0] zext_ln700_145_fu_11122_p1;
wire   [3:0] add_ln700_154_fu_11128_p2;
wire   [4:0] zext_ln700_149_fu_11134_p1;
wire   [4:0] zext_ln700_142_fu_11118_p1;
wire   [4:0] add_ln700_155_fu_11138_p2;
wire   [5:0] zext_ln700_150_fu_11144_p1;
wire   [5:0] zext_ln700_135_fu_11102_p1;
wire   [5:0] add_ln700_156_fu_11148_p2;
wire   [3:0] zext_ln700_157_fu_11161_p1;
wire   [3:0] zext_ln700_154_fu_11158_p1;
wire   [3:0] add_ln700_163_fu_11164_p2;
wire   [3:0] zext_ln700_164_fu_11177_p1;
wire   [3:0] zext_ln700_161_fu_11174_p1;
wire   [3:0] add_ln700_170_fu_11180_p2;
wire   [4:0] zext_ln700_165_fu_11186_p1;
wire   [4:0] zext_ln700_158_fu_11170_p1;
wire   [4:0] add_ln700_171_fu_11190_p2;
wire   [3:0] zext_ln700_172_fu_11203_p1;
wire   [3:0] zext_ln700_169_fu_11200_p1;
wire   [3:0] add_ln700_178_fu_11206_p2;
wire   [3:0] zext_ln700_179_fu_11219_p1;
wire   [3:0] zext_ln700_176_fu_11216_p1;
wire   [3:0] add_ln700_185_fu_11222_p2;
wire   [4:0] zext_ln700_180_fu_11228_p1;
wire   [4:0] zext_ln700_173_fu_11212_p1;
wire   [4:0] add_ln700_186_fu_11232_p2;
wire   [5:0] zext_ln700_181_fu_11238_p1;
wire   [5:0] zext_ln700_166_fu_11196_p1;
wire   [5:0] add_ln700_187_fu_11242_p2;
wire   [6:0] zext_ln700_182_fu_11248_p1;
wire   [6:0] zext_ln700_151_fu_11154_p1;
wire   [3:0] zext_ln700_189_fu_11261_p1;
wire   [3:0] zext_ln700_186_fu_11258_p1;
wire   [3:0] add_ln700_195_fu_11264_p2;
wire   [3:0] zext_ln700_196_fu_11277_p1;
wire   [3:0] zext_ln700_193_fu_11274_p1;
wire   [3:0] add_ln700_202_fu_11280_p2;
wire   [4:0] zext_ln700_197_fu_11286_p1;
wire   [4:0] zext_ln700_190_fu_11270_p1;
wire   [4:0] add_ln700_203_fu_11290_p2;
wire   [3:0] zext_ln700_204_fu_11303_p1;
wire   [3:0] zext_ln700_201_fu_11300_p1;
wire   [3:0] add_ln700_210_fu_11306_p2;
wire   [3:0] zext_ln700_211_fu_11319_p1;
wire   [3:0] zext_ln700_208_fu_11316_p1;
wire   [3:0] add_ln700_217_fu_11322_p2;
wire   [4:0] zext_ln700_212_fu_11328_p1;
wire   [4:0] zext_ln700_205_fu_11312_p1;
wire   [4:0] add_ln700_218_fu_11332_p2;
wire   [5:0] zext_ln700_213_fu_11338_p1;
wire   [5:0] zext_ln700_198_fu_11296_p1;
wire   [5:0] add_ln700_219_fu_11342_p2;
wire   [3:0] zext_ln700_220_fu_11355_p1;
wire   [3:0] zext_ln700_217_fu_11352_p1;
wire   [3:0] add_ln700_226_fu_11358_p2;
wire   [3:0] zext_ln700_227_fu_11371_p1;
wire   [3:0] zext_ln700_224_fu_11368_p1;
wire   [3:0] add_ln700_233_fu_11374_p2;
wire   [4:0] zext_ln700_228_fu_11380_p1;
wire   [4:0] zext_ln700_221_fu_11364_p1;
wire   [4:0] add_ln700_234_fu_11384_p2;
wire   [3:0] zext_ln700_235_fu_11397_p1;
wire   [3:0] zext_ln700_232_fu_11394_p1;
wire   [3:0] add_ln700_241_fu_11400_p2;
wire   [3:0] zext_ln700_242_fu_11413_p1;
wire   [3:0] zext_ln700_239_fu_11410_p1;
wire   [3:0] add_ln700_248_fu_11416_p2;
wire   [4:0] zext_ln700_243_fu_11422_p1;
wire   [4:0] zext_ln700_236_fu_11406_p1;
wire   [4:0] add_ln700_249_fu_11426_p2;
wire   [5:0] zext_ln700_244_fu_11432_p1;
wire   [5:0] zext_ln700_229_fu_11390_p1;
wire   [5:0] add_ln700_250_fu_11436_p2;
wire   [6:0] zext_ln700_245_fu_11442_p1;
wire   [6:0] zext_ln700_214_fu_11348_p1;
wire   [7:0] zext_ln700_26_fu_11452_p1;
wire   [7:0] zext_ln700_57_fu_11460_p1;
wire   [7:0] add_ln700_29_fu_11455_p2;
wire   [7:0] zext_ln700_120_fu_11469_p1;
wire   [7:0] add_ln700_61_fu_11463_p2;
wire   [7:0] zext_ln700_246_fu_11481_p1;
wire   [7:0] zext_ln700_183_fu_11478_p1;
wire   [7:0] add_ln700_252_fu_11484_p2;
wire   [7:0] add_ln700_125_fu_11472_p2;
wire    ap_CS_fsm_state6;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

Thresholding_Batch_0_Thresholding_Batcbkb #(
    .DataWidth( 1 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_254_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_254_address0),
    .ce0(threshs_m_thresholds_254_ce0),
    .q0(threshs_m_thresholds_254_q0)
);

Thresholding_Batch_0_Thresholding_Batccud #(
    .DataWidth( 2 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_253_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_253_address0),
    .ce0(threshs_m_thresholds_253_ce0),
    .q0(threshs_m_thresholds_253_q0)
);

Thresholding_Batch_0_Thresholding_Batcbkb #(
    .DataWidth( 1 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_142_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_142_address0),
    .ce0(threshs_m_thresholds_142_ce0),
    .q0(threshs_m_thresholds_142_q0)
);

Thresholding_Batch_0_Thresholding_BatceOg #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_76_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_76_address0),
    .ce0(threshs_m_thresholds_76_ce0),
    .q0(threshs_m_thresholds_76_q0)
);

Thresholding_Batch_0_Thresholding_BatcfYi #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_65_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_65_address0),
    .ce0(threshs_m_thresholds_65_ce0),
    .q0(threshs_m_thresholds_65_q0)
);

Thresholding_Batch_0_Thresholding_Batccud #(
    .DataWidth( 2 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_54_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_54_address0),
    .ce0(threshs_m_thresholds_54_ce0),
    .q0(threshs_m_thresholds_54_q0)
);

Thresholding_Batch_0_Thresholding_Batcbkb #(
    .DataWidth( 1 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_43_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_43_address0),
    .ce0(threshs_m_thresholds_43_ce0),
    .q0(threshs_m_thresholds_43_q0)
);

Thresholding_Batch_0_Thresholding_Batcibs #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_32_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_32_address0),
    .ce0(threshs_m_thresholds_32_ce0),
    .q0(threshs_m_thresholds_32_q0)
);

Thresholding_Batch_0_Thresholding_BatcjbC #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_21_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_21_address0),
    .ce0(threshs_m_thresholds_21_ce0),
    .q0(threshs_m_thresholds_21_q0)
);

Thresholding_Batch_0_Thresholding_BatckbM #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_10_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_10_address0),
    .ce0(threshs_m_thresholds_10_ce0),
    .q0(threshs_m_thresholds_10_q0)
);

Thresholding_Batch_0_Thresholding_BatclbW #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_252_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_252_address0),
    .ce0(threshs_m_thresholds_252_ce0),
    .q0(threshs_m_thresholds_252_q0)
);

Thresholding_Batch_0_Thresholding_BatceOg #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_241_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_241_address0),
    .ce0(threshs_m_thresholds_241_ce0),
    .q0(threshs_m_thresholds_241_q0)
);

Thresholding_Batch_0_Thresholding_BatcfYi #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_230_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_230_address0),
    .ce0(threshs_m_thresholds_230_ce0),
    .q0(threshs_m_thresholds_230_q0)
);

Thresholding_Batch_0_Thresholding_Batccud #(
    .DataWidth( 2 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_219_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_219_address0),
    .ce0(threshs_m_thresholds_219_ce0),
    .q0(threshs_m_thresholds_219_q0)
);

Thresholding_Batch_0_Thresholding_Batcbkb #(
    .DataWidth( 1 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_208_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_208_address0),
    .ce0(threshs_m_thresholds_208_ce0),
    .q0(threshs_m_thresholds_208_q0)
);

Thresholding_Batch_0_Thresholding_BatcqcK #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_197_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_197_address0),
    .ce0(threshs_m_thresholds_197_ce0),
    .q0(threshs_m_thresholds_197_q0)
);

Thresholding_Batch_0_Thresholding_BatcrcU #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_186_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_186_address0),
    .ce0(threshs_m_thresholds_186_ce0),
    .q0(threshs_m_thresholds_186_q0)
);

Thresholding_Batch_0_Thresholding_Batcsc4 #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_175_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_175_address0),
    .ce0(threshs_m_thresholds_175_ce0),
    .q0(threshs_m_thresholds_175_q0)
);

Thresholding_Batch_0_Thresholding_Batctde #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_164_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_164_address0),
    .ce0(threshs_m_thresholds_164_ce0),
    .q0(threshs_m_thresholds_164_q0)
);

Thresholding_Batch_0_Thresholding_Batcudo #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_153_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_153_address0),
    .ce0(threshs_m_thresholds_153_ce0),
    .q0(threshs_m_thresholds_153_q0)
);

Thresholding_Batch_0_Thresholding_Batcvdy #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_141_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_141_address0),
    .ce0(threshs_m_thresholds_141_ce0),
    .q0(threshs_m_thresholds_141_q0)
);

Thresholding_Batch_0_Thresholding_BatcwdI #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_130_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_130_address0),
    .ce0(threshs_m_thresholds_130_ce0),
    .q0(threshs_m_thresholds_130_q0)
);

Thresholding_Batch_0_Thresholding_BatcxdS #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_119_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_119_address0),
    .ce0(threshs_m_thresholds_119_ce0),
    .q0(threshs_m_thresholds_119_q0)
);

Thresholding_Batch_0_Thresholding_Batcibs #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_108_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_108_address0),
    .ce0(threshs_m_thresholds_108_ce0),
    .q0(threshs_m_thresholds_108_q0)
);

Thresholding_Batch_0_Thresholding_BatcjbC #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_97_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_97_address0),
    .ce0(threshs_m_thresholds_97_ce0),
    .q0(threshs_m_thresholds_97_q0)
);

Thresholding_Batch_0_Thresholding_BatckbM #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_86_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_86_address0),
    .ce0(threshs_m_thresholds_86_ce0),
    .q0(threshs_m_thresholds_86_q0)
);

Thresholding_Batch_0_Thresholding_BatclbW #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_80_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_80_address0),
    .ce0(threshs_m_thresholds_80_ce0),
    .q0(threshs_m_thresholds_80_q0)
);

Thresholding_Batch_0_Thresholding_BatceOg #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_79_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_79_address0),
    .ce0(threshs_m_thresholds_79_ce0),
    .q0(threshs_m_thresholds_79_q0)
);

Thresholding_Batch_0_Thresholding_BatcfYi #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_78_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_78_address0),
    .ce0(threshs_m_thresholds_78_ce0),
    .q0(threshs_m_thresholds_78_q0)
);

Thresholding_Batch_0_Thresholding_Batccud #(
    .DataWidth( 2 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_77_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_77_address0),
    .ce0(threshs_m_thresholds_77_ce0),
    .q0(threshs_m_thresholds_77_q0)
);

Thresholding_Batch_0_Thresholding_Batcbkb #(
    .DataWidth( 1 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_75_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_75_address0),
    .ce0(threshs_m_thresholds_75_ce0),
    .q0(threshs_m_thresholds_75_q0)
);

Thresholding_Batch_0_Thresholding_BatcGfk #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_74_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_74_address0),
    .ce0(threshs_m_thresholds_74_ce0),
    .q0(threshs_m_thresholds_74_q0)
);

Thresholding_Batch_0_Thresholding_BatcHfu #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_73_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_73_address0),
    .ce0(threshs_m_thresholds_73_ce0),
    .q0(threshs_m_thresholds_73_q0)
);

Thresholding_Batch_0_Thresholding_BatcIfE #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_72_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_72_address0),
    .ce0(threshs_m_thresholds_72_ce0),
    .q0(threshs_m_thresholds_72_q0)
);

Thresholding_Batch_0_Thresholding_BatcJfO #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_71_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_71_address0),
    .ce0(threshs_m_thresholds_71_ce0),
    .q0(threshs_m_thresholds_71_q0)
);

Thresholding_Batch_0_Thresholding_BatcKfY #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_70_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_70_address0),
    .ce0(threshs_m_thresholds_70_ce0),
    .q0(threshs_m_thresholds_70_q0)
);

Thresholding_Batch_0_Thresholding_BatcLf8 #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_69_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_69_address0),
    .ce0(threshs_m_thresholds_69_ce0),
    .q0(threshs_m_thresholds_69_q0)
);

Thresholding_Batch_0_Thresholding_BatcMgi #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_68_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_68_address0),
    .ce0(threshs_m_thresholds_68_ce0),
    .q0(threshs_m_thresholds_68_q0)
);

Thresholding_Batch_0_Thresholding_BatcNgs #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_67_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_67_address0),
    .ce0(threshs_m_thresholds_67_ce0),
    .q0(threshs_m_thresholds_67_q0)
);

Thresholding_Batch_0_Thresholding_BatcOgC #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_66_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_66_address0),
    .ce0(threshs_m_thresholds_66_ce0),
    .q0(threshs_m_thresholds_66_q0)
);

Thresholding_Batch_0_Thresholding_BatcPgM #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_64_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_64_address0),
    .ce0(threshs_m_thresholds_64_ce0),
    .q0(threshs_m_thresholds_64_q0)
);

Thresholding_Batch_0_Thresholding_BatcQgW #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_63_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_63_address0),
    .ce0(threshs_m_thresholds_63_ce0),
    .q0(threshs_m_thresholds_63_q0)
);

Thresholding_Batch_0_Thresholding_BatcRg6 #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_62_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_62_address0),
    .ce0(threshs_m_thresholds_62_ce0),
    .q0(threshs_m_thresholds_62_q0)
);

Thresholding_Batch_0_Thresholding_BatcShg #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_61_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_61_address0),
    .ce0(threshs_m_thresholds_61_ce0),
    .q0(threshs_m_thresholds_61_q0)
);

Thresholding_Batch_0_Thresholding_BatcThq #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_60_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_60_address0),
    .ce0(threshs_m_thresholds_60_ce0),
    .q0(threshs_m_thresholds_60_q0)
);

Thresholding_Batch_0_Thresholding_BatcUhA #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_59_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_59_address0),
    .ce0(threshs_m_thresholds_59_ce0),
    .q0(threshs_m_thresholds_59_q0)
);

Thresholding_Batch_0_Thresholding_BatcVhK #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_58_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_58_address0),
    .ce0(threshs_m_thresholds_58_ce0),
    .q0(threshs_m_thresholds_58_q0)
);

Thresholding_Batch_0_Thresholding_BatcqcK #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_57_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_57_address0),
    .ce0(threshs_m_thresholds_57_ce0),
    .q0(threshs_m_thresholds_57_q0)
);

Thresholding_Batch_0_Thresholding_BatcrcU #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_56_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_56_address0),
    .ce0(threshs_m_thresholds_56_ce0),
    .q0(threshs_m_thresholds_56_q0)
);

Thresholding_Batch_0_Thresholding_Batcsc4 #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_55_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_55_address0),
    .ce0(threshs_m_thresholds_55_ce0),
    .q0(threshs_m_thresholds_55_q0)
);

Thresholding_Batch_0_Thresholding_Batctde #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_53_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_53_address0),
    .ce0(threshs_m_thresholds_53_ce0),
    .q0(threshs_m_thresholds_53_q0)
);

Thresholding_Batch_0_Thresholding_Batcudo #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_52_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_52_address0),
    .ce0(threshs_m_thresholds_52_ce0),
    .q0(threshs_m_thresholds_52_q0)
);

Thresholding_Batch_0_Thresholding_Batcvdy #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_51_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_51_address0),
    .ce0(threshs_m_thresholds_51_ce0),
    .q0(threshs_m_thresholds_51_q0)
);

Thresholding_Batch_0_Thresholding_BatcwdI #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_50_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_50_address0),
    .ce0(threshs_m_thresholds_50_ce0),
    .q0(threshs_m_thresholds_50_q0)
);

Thresholding_Batch_0_Thresholding_BatcxdS #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_49_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_49_address0),
    .ce0(threshs_m_thresholds_49_ce0),
    .q0(threshs_m_thresholds_49_q0)
);

Thresholding_Batch_0_Thresholding_Batcibs #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_48_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_48_address0),
    .ce0(threshs_m_thresholds_48_ce0),
    .q0(threshs_m_thresholds_48_q0)
);

Thresholding_Batch_0_Thresholding_BatcjbC #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_47_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_47_address0),
    .ce0(threshs_m_thresholds_47_ce0),
    .q0(threshs_m_thresholds_47_q0)
);

Thresholding_Batch_0_Thresholding_BatckbM #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_46_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_46_address0),
    .ce0(threshs_m_thresholds_46_ce0),
    .q0(threshs_m_thresholds_46_q0)
);

Thresholding_Batch_0_Thresholding_BatclbW #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_45_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_45_address0),
    .ce0(threshs_m_thresholds_45_ce0),
    .q0(threshs_m_thresholds_45_q0)
);

Thresholding_Batch_0_Thresholding_BatceOg #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_44_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_44_address0),
    .ce0(threshs_m_thresholds_44_ce0),
    .q0(threshs_m_thresholds_44_q0)
);

Thresholding_Batch_0_Thresholding_BatcfYi #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_42_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_42_address0),
    .ce0(threshs_m_thresholds_42_ce0),
    .q0(threshs_m_thresholds_42_q0)
);

Thresholding_Batch_0_Thresholding_Batccud #(
    .DataWidth( 2 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_41_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_41_address0),
    .ce0(threshs_m_thresholds_41_ce0),
    .q0(threshs_m_thresholds_41_q0)
);

Thresholding_Batch_0_Thresholding_Batcbkb #(
    .DataWidth( 1 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_40_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_40_address0),
    .ce0(threshs_m_thresholds_40_ce0),
    .q0(threshs_m_thresholds_40_q0)
);

Thresholding_Batch_0_Thresholding_Batcbck #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_39_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_39_address0),
    .ce0(threshs_m_thresholds_39_ce0),
    .q0(threshs_m_thresholds_39_q0)
);

Thresholding_Batch_0_Thresholding_Batcbdk #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_38_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_38_address0),
    .ce0(threshs_m_thresholds_38_ce0),
    .q0(threshs_m_thresholds_38_q0)
);

Thresholding_Batch_0_Thresholding_Batcbek #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_37_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_37_address0),
    .ce0(threshs_m_thresholds_37_ce0),
    .q0(threshs_m_thresholds_37_q0)
);

Thresholding_Batch_0_Thresholding_Batcbfk #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_36_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_36_address0),
    .ce0(threshs_m_thresholds_36_ce0),
    .q0(threshs_m_thresholds_36_q0)
);

Thresholding_Batch_0_Thresholding_Batcbgk #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_35_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_35_address0),
    .ce0(threshs_m_thresholds_35_ce0),
    .q0(threshs_m_thresholds_35_q0)
);

Thresholding_Batch_0_Thresholding_Batcbhl #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_34_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_34_address0),
    .ce0(threshs_m_thresholds_34_ce0),
    .q0(threshs_m_thresholds_34_q0)
);

Thresholding_Batch_0_Thresholding_Batcbil #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_33_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_33_address0),
    .ce0(threshs_m_thresholds_33_ce0),
    .q0(threshs_m_thresholds_33_q0)
);

Thresholding_Batch_0_Thresholding_Batcbjl #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_31_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_31_address0),
    .ce0(threshs_m_thresholds_31_ce0),
    .q0(threshs_m_thresholds_31_q0)
);

Thresholding_Batch_0_Thresholding_Batcbkl #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_30_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_30_address0),
    .ce0(threshs_m_thresholds_30_ce0),
    .q0(threshs_m_thresholds_30_q0)
);

Thresholding_Batch_0_Thresholding_Batcbll #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_29_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_29_address0),
    .ce0(threshs_m_thresholds_29_ce0),
    .q0(threshs_m_thresholds_29_q0)
);

Thresholding_Batch_0_Thresholding_Batcbml #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_28_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_28_address0),
    .ce0(threshs_m_thresholds_28_ce0),
    .q0(threshs_m_thresholds_28_q0)
);

Thresholding_Batch_0_Thresholding_Batcbnm #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_27_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_27_address0),
    .ce0(threshs_m_thresholds_27_ce0),
    .q0(threshs_m_thresholds_27_q0)
);

Thresholding_Batch_0_Thresholding_Batcbom #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_26_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_26_address0),
    .ce0(threshs_m_thresholds_26_ce0),
    .q0(threshs_m_thresholds_26_q0)
);

Thresholding_Batch_0_Thresholding_Batcbpm #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_25_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_25_address0),
    .ce0(threshs_m_thresholds_25_ce0),
    .q0(threshs_m_thresholds_25_q0)
);

Thresholding_Batch_0_Thresholding_Batcbqm #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_24_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_24_address0),
    .ce0(threshs_m_thresholds_24_ce0),
    .q0(threshs_m_thresholds_24_q0)
);

Thresholding_Batch_0_Thresholding_Batcbrm #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_23_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_23_address0),
    .ce0(threshs_m_thresholds_23_ce0),
    .q0(threshs_m_thresholds_23_q0)
);

Thresholding_Batch_0_Thresholding_Batcbsm #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_22_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_22_address0),
    .ce0(threshs_m_thresholds_22_ce0),
    .q0(threshs_m_thresholds_22_q0)
);

Thresholding_Batch_0_Thresholding_Batcbtn #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_20_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_20_address0),
    .ce0(threshs_m_thresholds_20_ce0),
    .q0(threshs_m_thresholds_20_q0)
);

Thresholding_Batch_0_Thresholding_Batcbun #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_19_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_19_address0),
    .ce0(threshs_m_thresholds_19_ce0),
    .q0(threshs_m_thresholds_19_q0)
);

Thresholding_Batch_0_Thresholding_Batcbvn #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_18_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_18_address0),
    .ce0(threshs_m_thresholds_18_ce0),
    .q0(threshs_m_thresholds_18_q0)
);

Thresholding_Batch_0_Thresholding_Batcbwn #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_17_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_17_address0),
    .ce0(threshs_m_thresholds_17_ce0),
    .q0(threshs_m_thresholds_17_q0)
);

Thresholding_Batch_0_Thresholding_Batcbxn #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_16_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_16_address0),
    .ce0(threshs_m_thresholds_16_ce0),
    .q0(threshs_m_thresholds_16_q0)
);

Thresholding_Batch_0_Thresholding_Batcbyn #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_15_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_15_address0),
    .ce0(threshs_m_thresholds_15_ce0),
    .q0(threshs_m_thresholds_15_q0)
);

Thresholding_Batch_0_Thresholding_Batcbzo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_14_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_14_address0),
    .ce0(threshs_m_thresholds_14_ce0),
    .q0(threshs_m_thresholds_14_q0)
);

Thresholding_Batch_0_Thresholding_BatcbAo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_13_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_13_address0),
    .ce0(threshs_m_thresholds_13_ce0),
    .q0(threshs_m_thresholds_13_q0)
);

Thresholding_Batch_0_Thresholding_BatcbBo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_12_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_12_address0),
    .ce0(threshs_m_thresholds_12_ce0),
    .q0(threshs_m_thresholds_12_q0)
);

Thresholding_Batch_0_Thresholding_BatcbCo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_11_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_11_address0),
    .ce0(threshs_m_thresholds_11_ce0),
    .q0(threshs_m_thresholds_11_q0)
);

Thresholding_Batch_0_Thresholding_BatcbDo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_9_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_9_address0),
    .ce0(threshs_m_thresholds_9_ce0),
    .q0(threshs_m_thresholds_9_q0)
);

Thresholding_Batch_0_Thresholding_BatcbEo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_8_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_8_address0),
    .ce0(threshs_m_thresholds_8_ce0),
    .q0(threshs_m_thresholds_8_q0)
);

Thresholding_Batch_0_Thresholding_BatcbFp #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_7_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_7_address0),
    .ce0(threshs_m_thresholds_7_ce0),
    .q0(threshs_m_thresholds_7_q0)
);

Thresholding_Batch_0_Thresholding_BatcbGp #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_6_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_6_address0),
    .ce0(threshs_m_thresholds_6_ce0),
    .q0(threshs_m_thresholds_6_q0)
);

Thresholding_Batch_0_Thresholding_BatcbHp #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_5_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_5_address0),
    .ce0(threshs_m_thresholds_5_ce0),
    .q0(threshs_m_thresholds_5_q0)
);

Thresholding_Batch_0_Thresholding_BatcGfk #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_4_address0),
    .ce0(threshs_m_thresholds_4_ce0),
    .q0(threshs_m_thresholds_4_q0)
);

Thresholding_Batch_0_Thresholding_BatcHfu #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_3_address0),
    .ce0(threshs_m_thresholds_3_ce0),
    .q0(threshs_m_thresholds_3_q0)
);

Thresholding_Batch_0_Thresholding_BatcIfE #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_2_address0),
    .ce0(threshs_m_thresholds_2_ce0),
    .q0(threshs_m_thresholds_2_q0)
);

Thresholding_Batch_0_Thresholding_BatcJfO #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_1_address0),
    .ce0(threshs_m_thresholds_1_ce0),
    .q0(threshs_m_thresholds_1_q0)
);

Thresholding_Batch_0_Thresholding_BatcKfY #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_address0),
    .ce0(threshs_m_thresholds_ce0),
    .q0(threshs_m_thresholds_q0)
);

Thresholding_Batch_0_Thresholding_BatcLf8 #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_251_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_251_address0),
    .ce0(threshs_m_thresholds_251_ce0),
    .q0(threshs_m_thresholds_251_q0)
);

Thresholding_Batch_0_Thresholding_BatcMgi #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_250_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_250_address0),
    .ce0(threshs_m_thresholds_250_ce0),
    .q0(threshs_m_thresholds_250_q0)
);

Thresholding_Batch_0_Thresholding_BatcNgs #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_249_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_249_address0),
    .ce0(threshs_m_thresholds_249_ce0),
    .q0(threshs_m_thresholds_249_q0)
);

Thresholding_Batch_0_Thresholding_BatcOgC #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_248_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_248_address0),
    .ce0(threshs_m_thresholds_248_ce0),
    .q0(threshs_m_thresholds_248_q0)
);

Thresholding_Batch_0_Thresholding_BatcPgM #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_247_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_247_address0),
    .ce0(threshs_m_thresholds_247_ce0),
    .q0(threshs_m_thresholds_247_q0)
);

Thresholding_Batch_0_Thresholding_BatcQgW #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_246_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_246_address0),
    .ce0(threshs_m_thresholds_246_ce0),
    .q0(threshs_m_thresholds_246_q0)
);

Thresholding_Batch_0_Thresholding_BatcRg6 #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_245_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_245_address0),
    .ce0(threshs_m_thresholds_245_ce0),
    .q0(threshs_m_thresholds_245_q0)
);

Thresholding_Batch_0_Thresholding_BatcShg #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_244_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_244_address0),
    .ce0(threshs_m_thresholds_244_ce0),
    .q0(threshs_m_thresholds_244_q0)
);

Thresholding_Batch_0_Thresholding_BatcThq #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_243_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_243_address0),
    .ce0(threshs_m_thresholds_243_ce0),
    .q0(threshs_m_thresholds_243_q0)
);

Thresholding_Batch_0_Thresholding_BatcUhA #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_242_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_242_address0),
    .ce0(threshs_m_thresholds_242_ce0),
    .q0(threshs_m_thresholds_242_q0)
);

Thresholding_Batch_0_Thresholding_BatcVhK #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_240_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_240_address0),
    .ce0(threshs_m_thresholds_240_ce0),
    .q0(threshs_m_thresholds_240_q0)
);

Thresholding_Batch_0_Thresholding_BatcqcK #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_239_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_239_address0),
    .ce0(threshs_m_thresholds_239_ce0),
    .q0(threshs_m_thresholds_239_q0)
);

Thresholding_Batch_0_Thresholding_BatcrcU #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_238_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_238_address0),
    .ce0(threshs_m_thresholds_238_ce0),
    .q0(threshs_m_thresholds_238_q0)
);

Thresholding_Batch_0_Thresholding_Batcsc4 #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_237_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_237_address0),
    .ce0(threshs_m_thresholds_237_ce0),
    .q0(threshs_m_thresholds_237_q0)
);

Thresholding_Batch_0_Thresholding_Batctde #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_236_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_236_address0),
    .ce0(threshs_m_thresholds_236_ce0),
    .q0(threshs_m_thresholds_236_q0)
);

Thresholding_Batch_0_Thresholding_Batcudo #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_235_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_235_address0),
    .ce0(threshs_m_thresholds_235_ce0),
    .q0(threshs_m_thresholds_235_q0)
);

Thresholding_Batch_0_Thresholding_Batcvdy #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_234_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_234_address0),
    .ce0(threshs_m_thresholds_234_ce0),
    .q0(threshs_m_thresholds_234_q0)
);

Thresholding_Batch_0_Thresholding_BatcwdI #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_233_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_233_address0),
    .ce0(threshs_m_thresholds_233_ce0),
    .q0(threshs_m_thresholds_233_q0)
);

Thresholding_Batch_0_Thresholding_BatcxdS #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_232_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_232_address0),
    .ce0(threshs_m_thresholds_232_ce0),
    .q0(threshs_m_thresholds_232_q0)
);

Thresholding_Batch_0_Thresholding_Batcibs #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_231_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_231_address0),
    .ce0(threshs_m_thresholds_231_ce0),
    .q0(threshs_m_thresholds_231_q0)
);

Thresholding_Batch_0_Thresholding_BatcjbC #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_229_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_229_address0),
    .ce0(threshs_m_thresholds_229_ce0),
    .q0(threshs_m_thresholds_229_q0)
);

Thresholding_Batch_0_Thresholding_BatckbM #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_228_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_228_address0),
    .ce0(threshs_m_thresholds_228_ce0),
    .q0(threshs_m_thresholds_228_q0)
);

Thresholding_Batch_0_Thresholding_BatclbW #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_227_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_227_address0),
    .ce0(threshs_m_thresholds_227_ce0),
    .q0(threshs_m_thresholds_227_q0)
);

Thresholding_Batch_0_Thresholding_BatceOg #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_226_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_226_address0),
    .ce0(threshs_m_thresholds_226_ce0),
    .q0(threshs_m_thresholds_226_q0)
);

Thresholding_Batch_0_Thresholding_BatcfYi #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_225_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_225_address0),
    .ce0(threshs_m_thresholds_225_ce0),
    .q0(threshs_m_thresholds_225_q0)
);

Thresholding_Batch_0_Thresholding_Batccud #(
    .DataWidth( 2 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_224_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_224_address0),
    .ce0(threshs_m_thresholds_224_ce0),
    .q0(threshs_m_thresholds_224_q0)
);

Thresholding_Batch_0_Thresholding_Batcbkb #(
    .DataWidth( 1 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_223_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_223_address0),
    .ce0(threshs_m_thresholds_223_ce0),
    .q0(threshs_m_thresholds_223_q0)
);

Thresholding_Batch_0_Thresholding_Batcceu #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_222_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_222_address0),
    .ce0(threshs_m_thresholds_222_ce0),
    .q0(threshs_m_thresholds_222_q0)
);

Thresholding_Batch_0_Thresholding_Batcceu #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_221_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_221_address0),
    .ce0(threshs_m_thresholds_221_ce0),
    .q0(threshs_m_thresholds_221_q0)
);

Thresholding_Batch_0_Thresholding_Batccgu #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_220_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_220_address0),
    .ce0(threshs_m_thresholds_220_ce0),
    .q0(threshs_m_thresholds_220_q0)
);

Thresholding_Batch_0_Thresholding_Batcchv #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_218_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_218_address0),
    .ce0(threshs_m_thresholds_218_ce0),
    .q0(threshs_m_thresholds_218_q0)
);

Thresholding_Batch_0_Thresholding_Batcciv #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_217_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_217_address0),
    .ce0(threshs_m_thresholds_217_ce0),
    .q0(threshs_m_thresholds_217_q0)
);

Thresholding_Batch_0_Thresholding_Batccjv #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_216_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_216_address0),
    .ce0(threshs_m_thresholds_216_ce0),
    .q0(threshs_m_thresholds_216_q0)
);

Thresholding_Batch_0_Thresholding_Batcckv #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_215_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_215_address0),
    .ce0(threshs_m_thresholds_215_ce0),
    .q0(threshs_m_thresholds_215_q0)
);

Thresholding_Batch_0_Thresholding_Batcclv #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_214_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_214_address0),
    .ce0(threshs_m_thresholds_214_ce0),
    .q0(threshs_m_thresholds_214_q0)
);

Thresholding_Batch_0_Thresholding_Batccmv #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_213_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_213_address0),
    .ce0(threshs_m_thresholds_213_ce0),
    .q0(threshs_m_thresholds_213_q0)
);

Thresholding_Batch_0_Thresholding_Batccnw #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_212_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_212_address0),
    .ce0(threshs_m_thresholds_212_ce0),
    .q0(threshs_m_thresholds_212_q0)
);

Thresholding_Batch_0_Thresholding_Batccow #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_211_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_211_address0),
    .ce0(threshs_m_thresholds_211_ce0),
    .q0(threshs_m_thresholds_211_q0)
);

Thresholding_Batch_0_Thresholding_Batccpw #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_210_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_210_address0),
    .ce0(threshs_m_thresholds_210_ce0),
    .q0(threshs_m_thresholds_210_q0)
);

Thresholding_Batch_0_Thresholding_Batccqw #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_209_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_209_address0),
    .ce0(threshs_m_thresholds_209_ce0),
    .q0(threshs_m_thresholds_209_q0)
);

Thresholding_Batch_0_Thresholding_Batccrw #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_207_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_207_address0),
    .ce0(threshs_m_thresholds_207_ce0),
    .q0(threshs_m_thresholds_207_q0)
);

Thresholding_Batch_0_Thresholding_Batccsw #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_206_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_206_address0),
    .ce0(threshs_m_thresholds_206_ce0),
    .q0(threshs_m_thresholds_206_q0)
);

Thresholding_Batch_0_Thresholding_Batcctx #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_205_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_205_address0),
    .ce0(threshs_m_thresholds_205_ce0),
    .q0(threshs_m_thresholds_205_q0)
);

Thresholding_Batch_0_Thresholding_Batccux #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_204_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_204_address0),
    .ce0(threshs_m_thresholds_204_ce0),
    .q0(threshs_m_thresholds_204_q0)
);

Thresholding_Batch_0_Thresholding_Batccvx #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_203_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_203_address0),
    .ce0(threshs_m_thresholds_203_ce0),
    .q0(threshs_m_thresholds_203_q0)
);

Thresholding_Batch_0_Thresholding_Batccwx #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_202_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_202_address0),
    .ce0(threshs_m_thresholds_202_ce0),
    .q0(threshs_m_thresholds_202_q0)
);

Thresholding_Batch_0_Thresholding_Batccxx #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_201_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_201_address0),
    .ce0(threshs_m_thresholds_201_ce0),
    .q0(threshs_m_thresholds_201_q0)
);

Thresholding_Batch_0_Thresholding_Batccyx #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_200_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_200_address0),
    .ce0(threshs_m_thresholds_200_ce0),
    .q0(threshs_m_thresholds_200_q0)
);

Thresholding_Batch_0_Thresholding_Batcczy #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_199_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_199_address0),
    .ce0(threshs_m_thresholds_199_ce0),
    .q0(threshs_m_thresholds_199_q0)
);

Thresholding_Batch_0_Thresholding_BatccAy #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_198_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_198_address0),
    .ce0(threshs_m_thresholds_198_ce0),
    .q0(threshs_m_thresholds_198_q0)
);

Thresholding_Batch_0_Thresholding_BatccBy #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_196_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_196_address0),
    .ce0(threshs_m_thresholds_196_ce0),
    .q0(threshs_m_thresholds_196_q0)
);

Thresholding_Batch_0_Thresholding_BatccCy #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_195_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_195_address0),
    .ce0(threshs_m_thresholds_195_ce0),
    .q0(threshs_m_thresholds_195_q0)
);

Thresholding_Batch_0_Thresholding_BatccDy #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_194_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_194_address0),
    .ce0(threshs_m_thresholds_194_ce0),
    .q0(threshs_m_thresholds_194_q0)
);

Thresholding_Batch_0_Thresholding_BatccEy #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_193_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_193_address0),
    .ce0(threshs_m_thresholds_193_ce0),
    .q0(threshs_m_thresholds_193_q0)
);

Thresholding_Batch_0_Thresholding_BatccFz #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_192_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_192_address0),
    .ce0(threshs_m_thresholds_192_ce0),
    .q0(threshs_m_thresholds_192_q0)
);

Thresholding_Batch_0_Thresholding_BatccGz #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_191_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_191_address0),
    .ce0(threshs_m_thresholds_191_ce0),
    .q0(threshs_m_thresholds_191_q0)
);

Thresholding_Batch_0_Thresholding_BatccHz #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_190_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_190_address0),
    .ce0(threshs_m_thresholds_190_ce0),
    .q0(threshs_m_thresholds_190_q0)
);

Thresholding_Batch_0_Thresholding_BatccIz #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_189_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_189_address0),
    .ce0(threshs_m_thresholds_189_ce0),
    .q0(threshs_m_thresholds_189_q0)
);

Thresholding_Batch_0_Thresholding_BatccJz #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_188_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_188_address0),
    .ce0(threshs_m_thresholds_188_ce0),
    .q0(threshs_m_thresholds_188_q0)
);

Thresholding_Batch_0_Thresholding_BatccKz #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_187_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_187_address0),
    .ce0(threshs_m_thresholds_187_ce0),
    .q0(threshs_m_thresholds_187_q0)
);

Thresholding_Batch_0_Thresholding_BatccLz #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_185_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_185_address0),
    .ce0(threshs_m_thresholds_185_ce0),
    .q0(threshs_m_thresholds_185_q0)
);

Thresholding_Batch_0_Thresholding_BatccMA #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_184_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_184_address0),
    .ce0(threshs_m_thresholds_184_ce0),
    .q0(threshs_m_thresholds_184_q0)
);

Thresholding_Batch_0_Thresholding_BatccNA #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_183_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_183_address0),
    .ce0(threshs_m_thresholds_183_ce0),
    .q0(threshs_m_thresholds_183_q0)
);

Thresholding_Batch_0_Thresholding_BatccOA #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_182_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_182_address0),
    .ce0(threshs_m_thresholds_182_ce0),
    .q0(threshs_m_thresholds_182_q0)
);

Thresholding_Batch_0_Thresholding_BatccPA #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_181_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_181_address0),
    .ce0(threshs_m_thresholds_181_ce0),
    .q0(threshs_m_thresholds_181_q0)
);

Thresholding_Batch_0_Thresholding_BatccQA #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_180_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_180_address0),
    .ce0(threshs_m_thresholds_180_ce0),
    .q0(threshs_m_thresholds_180_q0)
);

Thresholding_Batch_0_Thresholding_BatccRA #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_179_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_179_address0),
    .ce0(threshs_m_thresholds_179_ce0),
    .q0(threshs_m_thresholds_179_q0)
);

Thresholding_Batch_0_Thresholding_BatccSB #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_178_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_178_address0),
    .ce0(threshs_m_thresholds_178_ce0),
    .q0(threshs_m_thresholds_178_q0)
);

Thresholding_Batch_0_Thresholding_BatccTB #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_177_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_177_address0),
    .ce0(threshs_m_thresholds_177_ce0),
    .q0(threshs_m_thresholds_177_q0)
);

Thresholding_Batch_0_Thresholding_BatccUB #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_176_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_176_address0),
    .ce0(threshs_m_thresholds_176_ce0),
    .q0(threshs_m_thresholds_176_q0)
);

Thresholding_Batch_0_Thresholding_BatccVB #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_174_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_174_address0),
    .ce0(threshs_m_thresholds_174_ce0),
    .q0(threshs_m_thresholds_174_q0)
);

Thresholding_Batch_0_Thresholding_BatccWB #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_173_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_173_address0),
    .ce0(threshs_m_thresholds_173_ce0),
    .q0(threshs_m_thresholds_173_q0)
);

Thresholding_Batch_0_Thresholding_BatccXB #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_172_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_172_address0),
    .ce0(threshs_m_thresholds_172_ce0),
    .q0(threshs_m_thresholds_172_q0)
);

Thresholding_Batch_0_Thresholding_BatccYC #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_171_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_171_address0),
    .ce0(threshs_m_thresholds_171_ce0),
    .q0(threshs_m_thresholds_171_q0)
);

Thresholding_Batch_0_Thresholding_BatccZC #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_170_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_170_address0),
    .ce0(threshs_m_thresholds_170_ce0),
    .q0(threshs_m_thresholds_170_q0)
);

Thresholding_Batch_0_Thresholding_Batcc0C #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_169_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_169_address0),
    .ce0(threshs_m_thresholds_169_ce0),
    .q0(threshs_m_thresholds_169_q0)
);

Thresholding_Batch_0_Thresholding_Batcc1C #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_168_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_168_address0),
    .ce0(threshs_m_thresholds_168_ce0),
    .q0(threshs_m_thresholds_168_q0)
);

Thresholding_Batch_0_Thresholding_Batcc2C #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_167_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_167_address0),
    .ce0(threshs_m_thresholds_167_ce0),
    .q0(threshs_m_thresholds_167_q0)
);

Thresholding_Batch_0_Thresholding_Batcc3C #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_166_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_166_address0),
    .ce0(threshs_m_thresholds_166_ce0),
    .q0(threshs_m_thresholds_166_q0)
);

Thresholding_Batch_0_Thresholding_Batcc4D #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_165_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_165_address0),
    .ce0(threshs_m_thresholds_165_ce0),
    .q0(threshs_m_thresholds_165_q0)
);

Thresholding_Batch_0_Thresholding_Batcc5D #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_163_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_163_address0),
    .ce0(threshs_m_thresholds_163_ce0),
    .q0(threshs_m_thresholds_163_q0)
);

Thresholding_Batch_0_Thresholding_Batcc6D #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_162_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_162_address0),
    .ce0(threshs_m_thresholds_162_ce0),
    .q0(threshs_m_thresholds_162_q0)
);

Thresholding_Batch_0_Thresholding_Batcc7D #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_161_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_161_address0),
    .ce0(threshs_m_thresholds_161_ce0),
    .q0(threshs_m_thresholds_161_q0)
);

Thresholding_Batch_0_Thresholding_Batcc8D #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_160_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_160_address0),
    .ce0(threshs_m_thresholds_160_ce0),
    .q0(threshs_m_thresholds_160_q0)
);

Thresholding_Batch_0_Thresholding_Batcc9D #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_159_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_159_address0),
    .ce0(threshs_m_thresholds_159_ce0),
    .q0(threshs_m_thresholds_159_q0)
);

Thresholding_Batch_0_Thresholding_BatcdaE #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_158_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_158_address0),
    .ce0(threshs_m_thresholds_158_ce0),
    .q0(threshs_m_thresholds_158_q0)
);

Thresholding_Batch_0_Thresholding_BatcdbE #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_157_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_157_address0),
    .ce0(threshs_m_thresholds_157_ce0),
    .q0(threshs_m_thresholds_157_q0)
);

Thresholding_Batch_0_Thresholding_BatcdcE #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_156_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_156_address0),
    .ce0(threshs_m_thresholds_156_ce0),
    .q0(threshs_m_thresholds_156_q0)
);

Thresholding_Batch_0_Thresholding_BatcddE #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_155_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_155_address0),
    .ce0(threshs_m_thresholds_155_ce0),
    .q0(threshs_m_thresholds_155_q0)
);

Thresholding_Batch_0_Thresholding_BatcdeE_x #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_154_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_154_address0),
    .ce0(threshs_m_thresholds_154_ce0),
    .q0(threshs_m_thresholds_154_q0)
);

Thresholding_Batch_0_Thresholding_BatcdfE #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_152_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_152_address0),
    .ce0(threshs_m_thresholds_152_ce0),
    .q0(threshs_m_thresholds_152_q0)
);

Thresholding_Batch_0_Thresholding_BatcdgE #(
    .DataWidth( 8 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_151_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_151_address0),
    .ce0(threshs_m_thresholds_151_ce0),
    .q0(threshs_m_thresholds_151_q0)
);

Thresholding_Batch_0_Thresholding_Batcbck #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_150_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_150_address0),
    .ce0(threshs_m_thresholds_150_ce0),
    .q0(threshs_m_thresholds_150_q0)
);

Thresholding_Batch_0_Thresholding_Batcbdk #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_149_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_149_address0),
    .ce0(threshs_m_thresholds_149_ce0),
    .q0(threshs_m_thresholds_149_q0)
);

Thresholding_Batch_0_Thresholding_Batcbek #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_148_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_148_address0),
    .ce0(threshs_m_thresholds_148_ce0),
    .q0(threshs_m_thresholds_148_q0)
);

Thresholding_Batch_0_Thresholding_Batcbfk #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_147_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_147_address0),
    .ce0(threshs_m_thresholds_147_ce0),
    .q0(threshs_m_thresholds_147_q0)
);

Thresholding_Batch_0_Thresholding_Batcbgk #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_146_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_146_address0),
    .ce0(threshs_m_thresholds_146_ce0),
    .q0(threshs_m_thresholds_146_q0)
);

Thresholding_Batch_0_Thresholding_Batcbhl #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_145_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_145_address0),
    .ce0(threshs_m_thresholds_145_ce0),
    .q0(threshs_m_thresholds_145_q0)
);

Thresholding_Batch_0_Thresholding_Batcbil #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_144_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_144_address0),
    .ce0(threshs_m_thresholds_144_ce0),
    .q0(threshs_m_thresholds_144_q0)
);

Thresholding_Batch_0_Thresholding_Batcbjl #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_143_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_143_address0),
    .ce0(threshs_m_thresholds_143_ce0),
    .q0(threshs_m_thresholds_143_q0)
);

Thresholding_Batch_0_Thresholding_Batcbkl #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_140_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_140_address0),
    .ce0(threshs_m_thresholds_140_ce0),
    .q0(threshs_m_thresholds_140_q0)
);

Thresholding_Batch_0_Thresholding_Batcbll #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_139_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_139_address0),
    .ce0(threshs_m_thresholds_139_ce0),
    .q0(threshs_m_thresholds_139_q0)
);

Thresholding_Batch_0_Thresholding_Batcbml #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_138_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_138_address0),
    .ce0(threshs_m_thresholds_138_ce0),
    .q0(threshs_m_thresholds_138_q0)
);

Thresholding_Batch_0_Thresholding_Batcbnm #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_137_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_137_address0),
    .ce0(threshs_m_thresholds_137_ce0),
    .q0(threshs_m_thresholds_137_q0)
);

Thresholding_Batch_0_Thresholding_Batcbom #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_136_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_136_address0),
    .ce0(threshs_m_thresholds_136_ce0),
    .q0(threshs_m_thresholds_136_q0)
);

Thresholding_Batch_0_Thresholding_Batcbpm #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_135_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_135_address0),
    .ce0(threshs_m_thresholds_135_ce0),
    .q0(threshs_m_thresholds_135_q0)
);

Thresholding_Batch_0_Thresholding_Batcbqm #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_134_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_134_address0),
    .ce0(threshs_m_thresholds_134_ce0),
    .q0(threshs_m_thresholds_134_q0)
);

Thresholding_Batch_0_Thresholding_Batcbrm #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_133_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_133_address0),
    .ce0(threshs_m_thresholds_133_ce0),
    .q0(threshs_m_thresholds_133_q0)
);

Thresholding_Batch_0_Thresholding_Batcbsm #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_132_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_132_address0),
    .ce0(threshs_m_thresholds_132_ce0),
    .q0(threshs_m_thresholds_132_q0)
);

Thresholding_Batch_0_Thresholding_Batcbtn #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_131_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_131_address0),
    .ce0(threshs_m_thresholds_131_ce0),
    .q0(threshs_m_thresholds_131_q0)
);

Thresholding_Batch_0_Thresholding_Batcbun #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_129_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_129_address0),
    .ce0(threshs_m_thresholds_129_ce0),
    .q0(threshs_m_thresholds_129_q0)
);

Thresholding_Batch_0_Thresholding_Batcbvn #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_128_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_128_address0),
    .ce0(threshs_m_thresholds_128_ce0),
    .q0(threshs_m_thresholds_128_q0)
);

Thresholding_Batch_0_Thresholding_Batcbwn #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_127_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_127_address0),
    .ce0(threshs_m_thresholds_127_ce0),
    .q0(threshs_m_thresholds_127_q0)
);

Thresholding_Batch_0_Thresholding_Batcbxn #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_126_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_126_address0),
    .ce0(threshs_m_thresholds_126_ce0),
    .q0(threshs_m_thresholds_126_q0)
);

Thresholding_Batch_0_Thresholding_Batcbyn #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_125_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_125_address0),
    .ce0(threshs_m_thresholds_125_ce0),
    .q0(threshs_m_thresholds_125_q0)
);

Thresholding_Batch_0_Thresholding_Batcbzo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_124_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_124_address0),
    .ce0(threshs_m_thresholds_124_ce0),
    .q0(threshs_m_thresholds_124_q0)
);

Thresholding_Batch_0_Thresholding_BatcbAo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_123_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_123_address0),
    .ce0(threshs_m_thresholds_123_ce0),
    .q0(threshs_m_thresholds_123_q0)
);

Thresholding_Batch_0_Thresholding_BatcbBo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_122_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_122_address0),
    .ce0(threshs_m_thresholds_122_ce0),
    .q0(threshs_m_thresholds_122_q0)
);

Thresholding_Batch_0_Thresholding_BatcbCo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_121_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_121_address0),
    .ce0(threshs_m_thresholds_121_ce0),
    .q0(threshs_m_thresholds_121_q0)
);

Thresholding_Batch_0_Thresholding_BatcbDo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_120_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_120_address0),
    .ce0(threshs_m_thresholds_120_ce0),
    .q0(threshs_m_thresholds_120_q0)
);

Thresholding_Batch_0_Thresholding_BatcbEo #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_118_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_118_address0),
    .ce0(threshs_m_thresholds_118_ce0),
    .q0(threshs_m_thresholds_118_q0)
);

Thresholding_Batch_0_Thresholding_BatcbFp #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_117_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_117_address0),
    .ce0(threshs_m_thresholds_117_ce0),
    .q0(threshs_m_thresholds_117_q0)
);

Thresholding_Batch_0_Thresholding_BatcbGp #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_116_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_116_address0),
    .ce0(threshs_m_thresholds_116_ce0),
    .q0(threshs_m_thresholds_116_q0)
);

Thresholding_Batch_0_Thresholding_BatcbHp #(
    .DataWidth( 7 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_115_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_115_address0),
    .ce0(threshs_m_thresholds_115_ce0),
    .q0(threshs_m_thresholds_115_q0)
);

Thresholding_Batch_0_Thresholding_BatcGfk #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_114_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_114_address0),
    .ce0(threshs_m_thresholds_114_ce0),
    .q0(threshs_m_thresholds_114_q0)
);

Thresholding_Batch_0_Thresholding_BatcHfu #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_113_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_113_address0),
    .ce0(threshs_m_thresholds_113_ce0),
    .q0(threshs_m_thresholds_113_q0)
);

Thresholding_Batch_0_Thresholding_BatcIfE #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_112_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_112_address0),
    .ce0(threshs_m_thresholds_112_ce0),
    .q0(threshs_m_thresholds_112_q0)
);

Thresholding_Batch_0_Thresholding_BatcJfO #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_111_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_111_address0),
    .ce0(threshs_m_thresholds_111_ce0),
    .q0(threshs_m_thresholds_111_q0)
);

Thresholding_Batch_0_Thresholding_BatcKfY #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_110_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_110_address0),
    .ce0(threshs_m_thresholds_110_ce0),
    .q0(threshs_m_thresholds_110_q0)
);

Thresholding_Batch_0_Thresholding_BatcLf8 #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_109_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_109_address0),
    .ce0(threshs_m_thresholds_109_ce0),
    .q0(threshs_m_thresholds_109_q0)
);

Thresholding_Batch_0_Thresholding_BatcMgi #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_107_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_107_address0),
    .ce0(threshs_m_thresholds_107_ce0),
    .q0(threshs_m_thresholds_107_q0)
);

Thresholding_Batch_0_Thresholding_BatcNgs #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_106_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_106_address0),
    .ce0(threshs_m_thresholds_106_ce0),
    .q0(threshs_m_thresholds_106_q0)
);

Thresholding_Batch_0_Thresholding_BatcOgC #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_105_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_105_address0),
    .ce0(threshs_m_thresholds_105_ce0),
    .q0(threshs_m_thresholds_105_q0)
);

Thresholding_Batch_0_Thresholding_BatcPgM #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_104_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_104_address0),
    .ce0(threshs_m_thresholds_104_ce0),
    .q0(threshs_m_thresholds_104_q0)
);

Thresholding_Batch_0_Thresholding_BatcQgW #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_103_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_103_address0),
    .ce0(threshs_m_thresholds_103_ce0),
    .q0(threshs_m_thresholds_103_q0)
);

Thresholding_Batch_0_Thresholding_BatcRg6 #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_102_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_102_address0),
    .ce0(threshs_m_thresholds_102_ce0),
    .q0(threshs_m_thresholds_102_q0)
);

Thresholding_Batch_0_Thresholding_BatcShg #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_101_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_101_address0),
    .ce0(threshs_m_thresholds_101_ce0),
    .q0(threshs_m_thresholds_101_q0)
);

Thresholding_Batch_0_Thresholding_BatcThq #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_100_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_100_address0),
    .ce0(threshs_m_thresholds_100_ce0),
    .q0(threshs_m_thresholds_100_q0)
);

Thresholding_Batch_0_Thresholding_BatcUhA #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_99_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_99_address0),
    .ce0(threshs_m_thresholds_99_ce0),
    .q0(threshs_m_thresholds_99_q0)
);

Thresholding_Batch_0_Thresholding_BatcVhK #(
    .DataWidth( 6 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_98_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_98_address0),
    .ce0(threshs_m_thresholds_98_ce0),
    .q0(threshs_m_thresholds_98_q0)
);

Thresholding_Batch_0_Thresholding_BatcqcK #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_96_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_96_address0),
    .ce0(threshs_m_thresholds_96_ce0),
    .q0(threshs_m_thresholds_96_q0)
);

Thresholding_Batch_0_Thresholding_BatcrcU #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_95_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_95_address0),
    .ce0(threshs_m_thresholds_95_ce0),
    .q0(threshs_m_thresholds_95_q0)
);

Thresholding_Batch_0_Thresholding_Batcsc4 #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_94_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_94_address0),
    .ce0(threshs_m_thresholds_94_ce0),
    .q0(threshs_m_thresholds_94_q0)
);

Thresholding_Batch_0_Thresholding_Batctde #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_93_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_93_address0),
    .ce0(threshs_m_thresholds_93_ce0),
    .q0(threshs_m_thresholds_93_q0)
);

Thresholding_Batch_0_Thresholding_Batcudo #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_92_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_92_address0),
    .ce0(threshs_m_thresholds_92_ce0),
    .q0(threshs_m_thresholds_92_q0)
);

Thresholding_Batch_0_Thresholding_Batcvdy #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_91_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_91_address0),
    .ce0(threshs_m_thresholds_91_ce0),
    .q0(threshs_m_thresholds_91_q0)
);

Thresholding_Batch_0_Thresholding_BatcwdI #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_90_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_90_address0),
    .ce0(threshs_m_thresholds_90_ce0),
    .q0(threshs_m_thresholds_90_q0)
);

Thresholding_Batch_0_Thresholding_BatcxdS #(
    .DataWidth( 5 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_89_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_89_address0),
    .ce0(threshs_m_thresholds_89_ce0),
    .q0(threshs_m_thresholds_89_q0)
);

Thresholding_Batch_0_Thresholding_Batcibs #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_88_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_88_address0),
    .ce0(threshs_m_thresholds_88_ce0),
    .q0(threshs_m_thresholds_88_q0)
);

Thresholding_Batch_0_Thresholding_BatcjbC #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_87_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_87_address0),
    .ce0(threshs_m_thresholds_87_ce0),
    .q0(threshs_m_thresholds_87_q0)
);

Thresholding_Batch_0_Thresholding_BatckbM #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_85_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_85_address0),
    .ce0(threshs_m_thresholds_85_ce0),
    .q0(threshs_m_thresholds_85_q0)
);

Thresholding_Batch_0_Thresholding_BatclbW #(
    .DataWidth( 4 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_84_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_84_address0),
    .ce0(threshs_m_thresholds_84_ce0),
    .q0(threshs_m_thresholds_84_q0)
);

Thresholding_Batch_0_Thresholding_BatceOg #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_83_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_83_address0),
    .ce0(threshs_m_thresholds_83_ce0),
    .q0(threshs_m_thresholds_83_q0)
);

Thresholding_Batch_0_Thresholding_BatcfYi #(
    .DataWidth( 3 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_82_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_82_address0),
    .ce0(threshs_m_thresholds_82_ce0),
    .q0(threshs_m_thresholds_82_q0)
);

Thresholding_Batch_0_Thresholding_Batccud #(
    .DataWidth( 2 ),
    .AddressRange( 3 ),
    .AddressWidth( 2 ))
threshs_m_thresholds_81_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_81_address0),
    .ce0(threshs_m_thresholds_81_ce0),
    .q0(threshs_m_thresholds_81_q0)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_3928_p2 == 1'd0))) begin
        i_0_reg_3917 <= i_fu_3934_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_reg_3917 <= 12'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_3928_p2 == 1'd0))) begin
        nf_assign_reg_3906 <= nf_1_fu_4211_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        nf_assign_reg_3906 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_reg_11497 == 1'd0))) begin
        add_ln700_102_reg_13185 <= add_ln700_102_fu_9696_p2;
        add_ln700_105_reg_13190 <= add_ln700_105_fu_9722_p2;
        add_ln700_110_reg_13195 <= add_ln700_110_fu_9748_p2;
        add_ln700_113_reg_13200 <= add_ln700_113_fu_9774_p2;
        add_ln700_117_reg_13205 <= add_ln700_117_fu_9800_p2;
        add_ln700_11_reg_13070 <= add_ln700_11_fu_9098_p2;
        add_ln700_120_reg_13210 <= add_ln700_120_fu_9826_p2;
        add_ln700_128_reg_13215 <= add_ln700_128_fu_9852_p2;
        add_ln700_131_reg_13220 <= add_ln700_131_fu_9878_p2;
        add_ln700_135_reg_13225 <= add_ln700_135_fu_9904_p2;
        add_ln700_138_reg_13230 <= add_ln700_138_fu_9930_p2;
        add_ln700_143_reg_13235 <= add_ln700_143_fu_9956_p2;
        add_ln700_146_reg_13240 <= add_ln700_146_fu_9982_p2;
        add_ln700_150_reg_13245 <= add_ln700_150_fu_10008_p2;
        add_ln700_153_reg_13250 <= add_ln700_153_fu_10034_p2;
        add_ln700_159_reg_13255 <= add_ln700_159_fu_10060_p2;
        add_ln700_162_reg_13260 <= add_ln700_162_fu_10086_p2;
        add_ln700_166_reg_13265 <= add_ln700_166_fu_10112_p2;
        add_ln700_169_reg_13270 <= add_ln700_169_fu_10138_p2;
        add_ln700_16_reg_13075 <= add_ln700_16_fu_9124_p2;
        add_ln700_174_reg_13275 <= add_ln700_174_fu_10164_p2;
        add_ln700_177_reg_13280 <= add_ln700_177_fu_10190_p2;
        add_ln700_181_reg_13285 <= add_ln700_181_fu_10216_p2;
        add_ln700_184_reg_13290 <= add_ln700_184_fu_10242_p2;
        add_ln700_191_reg_13295 <= add_ln700_191_fu_10268_p2;
        add_ln700_194_reg_13300 <= add_ln700_194_fu_10294_p2;
        add_ln700_198_reg_13305 <= add_ln700_198_fu_10320_p2;
        add_ln700_19_reg_13080 <= add_ln700_19_fu_9150_p2;
        add_ln700_201_reg_13310 <= add_ln700_201_fu_10346_p2;
        add_ln700_206_reg_13315 <= add_ln700_206_fu_10372_p2;
        add_ln700_209_reg_13320 <= add_ln700_209_fu_10398_p2;
        add_ln700_213_reg_13325 <= add_ln700_213_fu_10424_p2;
        add_ln700_216_reg_13330 <= add_ln700_216_fu_10450_p2;
        add_ln700_222_reg_13335 <= add_ln700_222_fu_10476_p2;
        add_ln700_225_reg_13340 <= add_ln700_225_fu_10502_p2;
        add_ln700_229_reg_13345 <= add_ln700_229_fu_10528_p2;
        add_ln700_232_reg_13350 <= add_ln700_232_fu_10554_p2;
        add_ln700_237_reg_13355 <= add_ln700_237_fu_10580_p2;
        add_ln700_23_reg_13085 <= add_ln700_23_fu_9176_p2;
        add_ln700_240_reg_13360 <= add_ln700_240_fu_10606_p2;
        add_ln700_244_reg_13365 <= add_ln700_244_fu_10632_p2;
        add_ln700_247_reg_13370 <= add_ln700_247_fu_10658_p2;
        add_ln700_26_reg_13090 <= add_ln700_26_fu_9202_p2;
        add_ln700_32_reg_13095 <= add_ln700_32_fu_9228_p2;
        add_ln700_35_reg_13100 <= add_ln700_35_fu_9254_p2;
        add_ln700_39_reg_13105 <= add_ln700_39_fu_9280_p2;
        add_ln700_42_reg_13110 <= add_ln700_42_fu_9306_p2;
        add_ln700_47_reg_13115 <= add_ln700_47_fu_9332_p2;
        add_ln700_4_reg_13060 <= add_ln700_4_fu_9046_p2;
        add_ln700_50_reg_13120 <= add_ln700_50_fu_9358_p2;
        add_ln700_54_reg_13125 <= add_ln700_54_fu_9384_p2;
        add_ln700_57_reg_13130 <= add_ln700_57_fu_9410_p2;
        add_ln700_64_reg_13135 <= add_ln700_64_fu_9436_p2;
        add_ln700_67_reg_13140 <= add_ln700_67_fu_9462_p2;
        add_ln700_71_reg_13145 <= add_ln700_71_fu_9488_p2;
        add_ln700_74_reg_13150 <= add_ln700_74_fu_9514_p2;
        add_ln700_79_reg_13155 <= add_ln700_79_fu_9540_p2;
        add_ln700_82_reg_13160 <= add_ln700_82_fu_9566_p2;
        add_ln700_86_reg_13165 <= add_ln700_86_fu_9592_p2;
        add_ln700_89_reg_13170 <= add_ln700_89_fu_9618_p2;
        add_ln700_8_reg_13065 <= add_ln700_8_fu_9072_p2;
        add_ln700_95_reg_13175 <= add_ln700_95_fu_9644_p2;
        add_ln700_98_reg_13180 <= add_ln700_98_fu_9670_p2;
        icmp_ln899_1_reg_13050 <= icmp_ln899_1_fu_4232_p2;
        icmp_ln899_2_reg_13055 <= icmp_ln899_2_fu_4245_p2;
        icmp_ln899_reg_13045 <= icmp_ln899_fu_4223_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_reg_11497_pp0_iter1_reg == 1'd0))) begin
        add_ln700_124_reg_13390 <= add_ln700_124_fu_11058_p2;
        add_ln700_13_reg_13375 <= add_ln700_13_fu_10736_p2;
        add_ln700_188_reg_13395 <= add_ln700_188_fu_11252_p2;
        add_ln700_251_reg_13400 <= add_ln700_251_fu_11446_p2;
        add_ln700_28_reg_13380 <= add_ln700_28_fu_10774_p2;
        add_ln700_60_reg_13385 <= add_ln700_60_fu_10864_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        icmp_ln221_reg_11497 <= icmp_ln221_fu_3928_p2;
        icmp_ln221_reg_11497_pp0_iter1_reg <= icmp_ln221_reg_11497;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln221_reg_11497_pp0_iter2_reg <= icmp_ln221_reg_11497_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_3928_p2 == 1'd0))) begin
        tmp_V_1_reg_11506 <= in_V_V_TDATA;
    end
end

always @ (*) begin
    if ((icmp_ln221_fu_3928_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state6) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln221_fu_3928_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_3928_p2 == 1'd0))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (icmp_ln221_reg_11497_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_reg_11497_pp0_iter2_reg == 1'd0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_100_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_100_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_101_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_101_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_102_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_102_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_103_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_103_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_104_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_104_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_105_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_105_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_106_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_106_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_107_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_107_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_108_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_108_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_109_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_109_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_10_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_10_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_110_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_110_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_111_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_111_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_112_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_112_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_113_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_113_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_114_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_114_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_115_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_115_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_116_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_116_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_117_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_117_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_118_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_118_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_119_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_119_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_11_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_11_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_120_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_120_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_121_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_121_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_122_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_122_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_123_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_123_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_124_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_124_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_125_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_125_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_126_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_126_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_127_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_127_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_128_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_128_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_129_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_129_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_12_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_12_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_130_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_130_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_131_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_131_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_132_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_132_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_133_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_133_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_134_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_134_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_135_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_135_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_136_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_136_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_137_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_137_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_138_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_138_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_139_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_139_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_13_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_13_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_140_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_140_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_141_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_141_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_142_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_142_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_143_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_143_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_144_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_144_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_145_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_145_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_146_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_146_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_147_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_147_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_148_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_148_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_149_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_149_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_14_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_14_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_150_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_150_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_151_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_151_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_152_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_152_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_153_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_153_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_154_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_154_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_155_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_155_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_156_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_156_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_157_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_157_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_158_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_158_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_159_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_159_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_15_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_15_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_160_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_160_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_161_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_161_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_162_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_162_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_163_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_163_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_164_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_164_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_165_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_165_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_166_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_166_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_167_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_167_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_168_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_168_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_169_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_169_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_16_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_16_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_170_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_170_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_171_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_171_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_172_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_172_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_173_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_173_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_174_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_174_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_175_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_175_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_176_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_176_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_177_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_177_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_178_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_178_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_179_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_179_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_17_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_17_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_180_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_180_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_181_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_181_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_182_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_182_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_183_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_183_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_184_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_184_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_185_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_185_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_186_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_186_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_187_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_187_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_188_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_188_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_189_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_189_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_18_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_18_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_190_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_190_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_191_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_191_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_192_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_192_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_193_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_193_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_194_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_194_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_195_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_195_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_196_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_196_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_197_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_197_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_198_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_198_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_199_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_199_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_19_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_19_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_1_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_1_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_200_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_200_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_201_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_201_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_202_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_202_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_203_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_203_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_204_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_204_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_205_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_205_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_206_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_206_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_207_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_207_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_208_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_208_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_209_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_209_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_20_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_20_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_210_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_210_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_211_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_211_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_212_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_212_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_213_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_213_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_214_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_214_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_215_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_215_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_216_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_216_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_217_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_217_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_218_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_218_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_219_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_219_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_21_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_21_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_220_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_220_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_221_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_221_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_222_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_222_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_223_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_223_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_224_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_224_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_225_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_225_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_226_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_226_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_227_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_227_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_228_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_228_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_229_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_229_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_22_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_22_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_230_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_230_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_231_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_231_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_232_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_232_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_233_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_233_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_234_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_234_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_235_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_235_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_236_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_236_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_237_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_237_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_238_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_238_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_239_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_239_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_23_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_23_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_240_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_240_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_241_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_241_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_242_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_242_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_243_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_243_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_244_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_244_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_245_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_245_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_246_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_246_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_247_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_247_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_248_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_248_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_249_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_249_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_24_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_24_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_250_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_250_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_251_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_251_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_252_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_252_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_253_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_253_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_254_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_254_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_25_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_25_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_26_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_26_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_27_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_27_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_28_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_28_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_29_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_29_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_2_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_2_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_30_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_30_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_31_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_31_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_32_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_32_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_33_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_33_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_34_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_34_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_35_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_35_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_36_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_36_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_37_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_37_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_38_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_38_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_39_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_39_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_3_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_3_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_40_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_40_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_41_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_41_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_42_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_42_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_43_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_43_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_44_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_44_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_45_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_45_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_46_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_46_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_47_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_47_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_48_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_48_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_49_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_49_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_4_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_4_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_50_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_50_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_51_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_51_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_52_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_52_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_53_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_53_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_54_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_54_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_55_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_55_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_56_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_56_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_57_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_57_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_58_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_58_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_59_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_59_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_5_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_5_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_60_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_60_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_61_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_61_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_62_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_62_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_63_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_63_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_64_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_64_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_65_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_65_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_66_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_66_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_67_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_67_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_68_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_68_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_69_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_69_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_6_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_6_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_70_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_70_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_71_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_71_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_72_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_72_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_73_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_73_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_74_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_74_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_75_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_75_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_76_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_76_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_77_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_77_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_78_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_78_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_79_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_79_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_7_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_7_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_80_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_80_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_81_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_81_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_82_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_82_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_83_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_83_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_84_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_84_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_85_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_85_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_86_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_86_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_87_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_87_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_88_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_88_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_89_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_89_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_8_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_8_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_90_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_90_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_91_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_91_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_92_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_92_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_93_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_93_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_94_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_94_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_95_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_95_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_96_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_96_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_97_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_97_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_98_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_98_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_99_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_99_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_9_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_9_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_3928_p2 == 1'd1)) & ~((ap_enable_reg_pp0_iter2 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter2 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_3928_p2 == 1'd1)))) begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln700_100_fu_9676_p2 = (zext_ln142_202_fu_6321_p1 + zext_ln142_204_fu_6344_p1);

assign add_ln700_101_fu_9686_p2 = (zext_ln142_206_fu_6367_p1 + zext_ln142_208_fu_6390_p1);

assign add_ln700_102_fu_9696_p2 = (zext_ln700_97_fu_9692_p1 + zext_ln700_96_fu_9682_p1);

assign add_ln700_103_fu_9702_p2 = (zext_ln142_210_fu_6413_p1 + zext_ln142_212_fu_6436_p1);

assign add_ln700_104_fu_9712_p2 = (zext_ln142_214_fu_6459_p1 + zext_ln142_216_fu_6482_p1);

assign add_ln700_105_fu_9722_p2 = (zext_ln700_100_fu_9718_p1 + zext_ln700_99_fu_9708_p1);

assign add_ln700_106_fu_10986_p2 = (zext_ln700_101_fu_10983_p1 + zext_ln700_98_fu_10980_p1);

assign add_ln700_107_fu_10996_p2 = (zext_ln700_102_fu_10992_p1 + zext_ln700_95_fu_10976_p1);

assign add_ln700_108_fu_9728_p2 = (zext_ln142_218_fu_6505_p1 + zext_ln142_220_fu_6528_p1);

assign add_ln700_109_fu_9738_p2 = (zext_ln142_222_fu_6551_p1 + zext_ln142_224_fu_6574_p1);

assign add_ln700_10_fu_9088_p2 = (zext_ln142_25_fu_4475_p1 + zext_ln142_26_fu_4498_p1);

assign add_ln700_110_fu_9748_p2 = (zext_ln700_105_fu_9744_p1 + zext_ln700_104_fu_9734_p1);

assign add_ln700_111_fu_9754_p2 = (zext_ln142_226_fu_6597_p1 + zext_ln142_228_fu_6620_p1);

assign add_ln700_112_fu_9764_p2 = (zext_ln142_230_fu_6643_p1 + zext_ln142_232_fu_6666_p1);

assign add_ln700_113_fu_9774_p2 = (zext_ln700_108_fu_9770_p1 + zext_ln700_107_fu_9760_p1);

assign add_ln700_114_fu_11012_p2 = (zext_ln700_109_fu_11009_p1 + zext_ln700_106_fu_11006_p1);

assign add_ln700_115_fu_9780_p2 = (zext_ln142_234_fu_6689_p1 + zext_ln142_236_fu_6712_p1);

assign add_ln700_116_fu_9790_p2 = (zext_ln142_238_fu_6735_p1 + zext_ln142_240_fu_6758_p1);

assign add_ln700_117_fu_9800_p2 = (zext_ln700_112_fu_9796_p1 + zext_ln700_111_fu_9786_p1);

assign add_ln700_118_fu_9806_p2 = (zext_ln142_242_fu_6781_p1 + zext_ln142_244_fu_6804_p1);

assign add_ln700_119_fu_9816_p2 = (zext_ln142_246_fu_6827_p1 + zext_ln142_247_fu_6850_p1);

assign add_ln700_11_fu_9098_p2 = (zext_ln700_9_fu_9094_p1 + zext_ln700_8_fu_9084_p1);

assign add_ln700_120_fu_9826_p2 = (zext_ln700_115_fu_9822_p1 + zext_ln700_114_fu_9812_p1);

assign add_ln700_121_fu_11028_p2 = (zext_ln700_116_fu_11025_p1 + zext_ln700_113_fu_11022_p1);

assign add_ln700_122_fu_11038_p2 = (zext_ln700_117_fu_11034_p1 + zext_ln700_110_fu_11018_p1);

assign add_ln700_123_fu_11048_p2 = (zext_ln700_118_fu_11044_p1 + zext_ln700_103_fu_11002_p1);

assign add_ln700_124_fu_11058_p2 = (zext_ln700_119_fu_11054_p1 + zext_ln700_88_fu_10960_p1);

assign add_ln700_125_fu_11472_p2 = (zext_ln700_120_fu_11469_p1 + add_ln700_61_fu_11463_p2);

assign add_ln700_126_fu_9832_p2 = (zext_ln142_248_fu_6865_p1 + zext_ln142_249_fu_6880_p1);

assign add_ln700_127_fu_9842_p2 = (zext_ln142_250_fu_6895_p1 + zext_ln142_251_fu_6910_p1);

assign add_ln700_128_fu_9852_p2 = (zext_ln700_122_fu_9848_p1 + zext_ln700_121_fu_9838_p1);

assign add_ln700_129_fu_9858_p2 = (zext_ln142_252_fu_6925_p1 + zext_ln142_253_fu_6940_p1);

assign add_ln700_12_fu_10726_p2 = (zext_ln700_10_fu_10723_p1 + zext_ln700_7_fu_10720_p1);

assign add_ln700_130_fu_9868_p2 = (zext_ln142_254_fu_6955_p1 + zext_ln142_255_fu_6970_p1);

assign add_ln700_131_fu_9878_p2 = (zext_ln700_125_fu_9874_p1 + zext_ln700_124_fu_9864_p1);

assign add_ln700_132_fu_11070_p2 = (zext_ln700_126_fu_11067_p1 + zext_ln700_123_fu_11064_p1);

assign add_ln700_133_fu_9884_p2 = (zext_ln142_256_fu_6985_p1 + zext_ln142_257_fu_7000_p1);

assign add_ln700_134_fu_9894_p2 = (zext_ln142_258_fu_7015_p1 + zext_ln142_259_fu_7030_p1);

assign add_ln700_135_fu_9904_p2 = (zext_ln700_129_fu_9900_p1 + zext_ln700_128_fu_9890_p1);

assign add_ln700_136_fu_9910_p2 = (zext_ln142_260_fu_7045_p1 + zext_ln142_261_fu_7060_p1);

assign add_ln700_137_fu_9920_p2 = (zext_ln142_262_fu_7075_p1 + zext_ln142_263_fu_7090_p1);

assign add_ln700_138_fu_9930_p2 = (zext_ln700_132_fu_9926_p1 + zext_ln700_131_fu_9916_p1);

assign add_ln700_139_fu_11086_p2 = (zext_ln700_133_fu_11083_p1 + zext_ln700_130_fu_11080_p1);

assign add_ln700_13_fu_10736_p2 = (zext_ln700_11_fu_10732_p1 + add_ln700_5_fu_10714_p2);

assign add_ln700_140_fu_11096_p2 = (zext_ln700_134_fu_11092_p1 + zext_ln700_127_fu_11076_p1);

assign add_ln700_141_fu_9936_p2 = (zext_ln142_264_fu_7105_p1 + zext_ln142_265_fu_7120_p1);

assign add_ln700_142_fu_9946_p2 = (zext_ln142_266_fu_7135_p1 + zext_ln142_267_fu_7150_p1);

assign add_ln700_143_fu_9956_p2 = (zext_ln700_137_fu_9952_p1 + zext_ln700_136_fu_9942_p1);

assign add_ln700_144_fu_9962_p2 = (zext_ln142_268_fu_7165_p1 + zext_ln142_269_fu_7180_p1);

assign add_ln700_145_fu_9972_p2 = (zext_ln142_270_fu_7195_p1 + zext_ln142_271_fu_7210_p1);

assign add_ln700_146_fu_9982_p2 = (zext_ln700_140_fu_9978_p1 + zext_ln700_139_fu_9968_p1);

assign add_ln700_147_fu_11112_p2 = (zext_ln700_141_fu_11109_p1 + zext_ln700_138_fu_11106_p1);

assign add_ln700_148_fu_9988_p2 = (zext_ln142_272_fu_7225_p1 + zext_ln142_273_fu_7240_p1);

assign add_ln700_149_fu_9998_p2 = (zext_ln142_274_fu_7255_p1 + zext_ln142_275_fu_7270_p1);

assign add_ln700_14_fu_9104_p2 = (zext_ln142_28_fu_4517_p1 + zext_ln142_30_fu_4536_p1);

assign add_ln700_150_fu_10008_p2 = (zext_ln700_144_fu_10004_p1 + zext_ln700_143_fu_9994_p1);

assign add_ln700_151_fu_10014_p2 = (zext_ln142_276_fu_7285_p1 + zext_ln142_277_fu_7300_p1);

assign add_ln700_152_fu_10024_p2 = (zext_ln142_278_fu_7315_p1 + zext_ln142_279_fu_7330_p1);

assign add_ln700_153_fu_10034_p2 = (zext_ln700_147_fu_10030_p1 + zext_ln700_146_fu_10020_p1);

assign add_ln700_154_fu_11128_p2 = (zext_ln700_148_fu_11125_p1 + zext_ln700_145_fu_11122_p1);

assign add_ln700_155_fu_11138_p2 = (zext_ln700_149_fu_11134_p1 + zext_ln700_142_fu_11118_p1);

assign add_ln700_156_fu_11148_p2 = (zext_ln700_150_fu_11144_p1 + zext_ln700_135_fu_11102_p1);

assign add_ln700_157_fu_10040_p2 = (zext_ln142_280_fu_7345_p1 + zext_ln142_281_fu_7360_p1);

assign add_ln700_158_fu_10050_p2 = (zext_ln142_282_fu_7375_p1 + zext_ln142_283_fu_7390_p1);

assign add_ln700_159_fu_10060_p2 = (zext_ln700_153_fu_10056_p1 + zext_ln700_152_fu_10046_p1);

assign add_ln700_15_fu_9114_p2 = (zext_ln142_32_fu_4555_p1 + zext_ln142_34_fu_4574_p1);

assign add_ln700_160_fu_10066_p2 = (zext_ln142_284_fu_7405_p1 + zext_ln142_285_fu_7420_p1);

assign add_ln700_161_fu_10076_p2 = (zext_ln142_286_fu_7435_p1 + zext_ln142_287_fu_7450_p1);

assign add_ln700_162_fu_10086_p2 = (zext_ln700_156_fu_10082_p1 + zext_ln700_155_fu_10072_p1);

assign add_ln700_163_fu_11164_p2 = (zext_ln700_157_fu_11161_p1 + zext_ln700_154_fu_11158_p1);

assign add_ln700_164_fu_10092_p2 = (zext_ln142_288_fu_7465_p1 + zext_ln142_289_fu_7480_p1);

assign add_ln700_165_fu_10102_p2 = (zext_ln142_290_fu_7495_p1 + zext_ln142_291_fu_7510_p1);

assign add_ln700_166_fu_10112_p2 = (zext_ln700_160_fu_10108_p1 + zext_ln700_159_fu_10098_p1);

assign add_ln700_167_fu_10118_p2 = (zext_ln142_292_fu_7525_p1 + zext_ln142_293_fu_7540_p1);

assign add_ln700_168_fu_10128_p2 = (zext_ln142_294_fu_7555_p1 + zext_ln142_295_fu_7570_p1);

assign add_ln700_169_fu_10138_p2 = (zext_ln700_163_fu_10134_p1 + zext_ln700_162_fu_10124_p1);

assign add_ln700_16_fu_9124_p2 = (zext_ln700_13_fu_9120_p1 + zext_ln700_12_fu_9110_p1);

assign add_ln700_170_fu_11180_p2 = (zext_ln700_164_fu_11177_p1 + zext_ln700_161_fu_11174_p1);

assign add_ln700_171_fu_11190_p2 = (zext_ln700_165_fu_11186_p1 + zext_ln700_158_fu_11170_p1);

assign add_ln700_172_fu_10144_p2 = (zext_ln142_296_fu_7585_p1 + zext_ln142_297_fu_7600_p1);

assign add_ln700_173_fu_10154_p2 = (zext_ln142_298_fu_7615_p1 + zext_ln142_299_fu_7630_p1);

assign add_ln700_174_fu_10164_p2 = (zext_ln700_168_fu_10160_p1 + zext_ln700_167_fu_10150_p1);

assign add_ln700_175_fu_10170_p2 = (zext_ln142_300_fu_7645_p1 + zext_ln142_301_fu_7660_p1);

assign add_ln700_176_fu_10180_p2 = (zext_ln142_302_fu_7675_p1 + zext_ln142_303_fu_7690_p1);

assign add_ln700_177_fu_10190_p2 = (zext_ln700_171_fu_10186_p1 + zext_ln700_170_fu_10176_p1);

assign add_ln700_178_fu_11206_p2 = (zext_ln700_172_fu_11203_p1 + zext_ln700_169_fu_11200_p1);

assign add_ln700_179_fu_10196_p2 = (zext_ln142_304_fu_7705_p1 + zext_ln142_305_fu_7720_p1);

assign add_ln700_17_fu_9130_p2 = (zext_ln142_36_fu_4593_p1 + zext_ln142_38_fu_4612_p1);

assign add_ln700_180_fu_10206_p2 = (zext_ln142_306_fu_7735_p1 + zext_ln142_307_fu_7750_p1);

assign add_ln700_181_fu_10216_p2 = (zext_ln700_175_fu_10212_p1 + zext_ln700_174_fu_10202_p1);

assign add_ln700_182_fu_10222_p2 = (zext_ln142_308_fu_7765_p1 + zext_ln142_309_fu_7780_p1);

assign add_ln700_183_fu_10232_p2 = (zext_ln142_310_fu_7795_p1 + zext_ln142_311_fu_7810_p1);

assign add_ln700_184_fu_10242_p2 = (zext_ln700_178_fu_10238_p1 + zext_ln700_177_fu_10228_p1);

assign add_ln700_185_fu_11222_p2 = (zext_ln700_179_fu_11219_p1 + zext_ln700_176_fu_11216_p1);

assign add_ln700_186_fu_11232_p2 = (zext_ln700_180_fu_11228_p1 + zext_ln700_173_fu_11212_p1);

assign add_ln700_187_fu_11242_p2 = (zext_ln700_181_fu_11238_p1 + zext_ln700_166_fu_11196_p1);

assign add_ln700_188_fu_11252_p2 = (zext_ln700_182_fu_11248_p1 + zext_ln700_151_fu_11154_p1);

assign add_ln700_189_fu_10248_p2 = (zext_ln142_312_fu_7825_p1 + zext_ln142_313_fu_7844_p1);

assign add_ln700_18_fu_9140_p2 = (zext_ln142_40_fu_4631_p1 + zext_ln142_42_fu_4650_p1);

assign add_ln700_190_fu_10258_p2 = (zext_ln142_314_fu_7863_p1 + zext_ln142_315_fu_7882_p1);

assign add_ln700_191_fu_10268_p2 = (zext_ln700_185_fu_10264_p1 + zext_ln700_184_fu_10254_p1);

assign add_ln700_192_fu_10274_p2 = (zext_ln142_316_fu_7901_p1 + zext_ln142_317_fu_7920_p1);

assign add_ln700_193_fu_10284_p2 = (zext_ln142_318_fu_7939_p1 + zext_ln142_319_fu_7958_p1);

assign add_ln700_194_fu_10294_p2 = (zext_ln700_188_fu_10290_p1 + zext_ln700_187_fu_10280_p1);

assign add_ln700_195_fu_11264_p2 = (zext_ln700_189_fu_11261_p1 + zext_ln700_186_fu_11258_p1);

assign add_ln700_196_fu_10300_p2 = (zext_ln142_320_fu_7977_p1 + zext_ln142_321_fu_7996_p1);

assign add_ln700_197_fu_10310_p2 = (zext_ln142_322_fu_8015_p1 + zext_ln142_323_fu_8034_p1);

assign add_ln700_198_fu_10320_p2 = (zext_ln700_192_fu_10316_p1 + zext_ln700_191_fu_10306_p1);

assign add_ln700_199_fu_10326_p2 = (zext_ln142_324_fu_8053_p1 + zext_ln142_325_fu_8072_p1);

assign add_ln700_19_fu_9150_p2 = (zext_ln700_16_fu_9146_p1 + zext_ln700_15_fu_9136_p1);

assign add_ln700_1_fu_10705_p2 = (zext_ln700_1_fu_10701_p1 + or_ln_fu_10669_p3);

assign add_ln700_200_fu_10336_p2 = (zext_ln142_326_fu_8091_p1 + zext_ln142_327_fu_8110_p1);

assign add_ln700_201_fu_10346_p2 = (zext_ln700_195_fu_10342_p1 + zext_ln700_194_fu_10332_p1);

assign add_ln700_202_fu_11280_p2 = (zext_ln700_196_fu_11277_p1 + zext_ln700_193_fu_11274_p1);

assign add_ln700_203_fu_11290_p2 = (zext_ln700_197_fu_11286_p1 + zext_ln700_190_fu_11270_p1);

assign add_ln700_204_fu_10352_p2 = (zext_ln142_328_fu_8129_p1 + zext_ln142_329_fu_8148_p1);

assign add_ln700_205_fu_10362_p2 = (zext_ln142_330_fu_8167_p1 + zext_ln142_331_fu_8186_p1);

assign add_ln700_206_fu_10372_p2 = (zext_ln700_200_fu_10368_p1 + zext_ln700_199_fu_10358_p1);

assign add_ln700_207_fu_10378_p2 = (zext_ln142_332_fu_8205_p1 + zext_ln142_333_fu_8224_p1);

assign add_ln700_208_fu_10388_p2 = (zext_ln142_334_fu_8243_p1 + zext_ln142_335_fu_8262_p1);

assign add_ln700_209_fu_10398_p2 = (zext_ln700_203_fu_10394_p1 + zext_ln700_202_fu_10384_p1);

assign add_ln700_20_fu_10748_p2 = (zext_ln700_17_fu_10745_p1 + zext_ln700_14_fu_10742_p1);

assign add_ln700_210_fu_11306_p2 = (zext_ln700_204_fu_11303_p1 + zext_ln700_201_fu_11300_p1);

assign add_ln700_211_fu_10404_p2 = (zext_ln142_336_fu_8281_p1 + zext_ln142_337_fu_8300_p1);

assign add_ln700_212_fu_10414_p2 = (zext_ln142_338_fu_8319_p1 + zext_ln142_339_fu_8338_p1);

assign add_ln700_213_fu_10424_p2 = (zext_ln700_207_fu_10420_p1 + zext_ln700_206_fu_10410_p1);

assign add_ln700_214_fu_10430_p2 = (zext_ln142_340_fu_8357_p1 + zext_ln142_341_fu_8376_p1);

assign add_ln700_215_fu_10440_p2 = (zext_ln142_342_fu_8395_p1 + zext_ln142_343_fu_8414_p1);

assign add_ln700_216_fu_10450_p2 = (zext_ln700_210_fu_10446_p1 + zext_ln700_209_fu_10436_p1);

assign add_ln700_217_fu_11322_p2 = (zext_ln700_211_fu_11319_p1 + zext_ln700_208_fu_11316_p1);

assign add_ln700_218_fu_11332_p2 = (zext_ln700_212_fu_11328_p1 + zext_ln700_205_fu_11312_p1);

assign add_ln700_219_fu_11342_p2 = (zext_ln700_213_fu_11338_p1 + zext_ln700_198_fu_11296_p1);

assign add_ln700_21_fu_9156_p2 = (zext_ln142_44_fu_4673_p1 + zext_ln142_46_fu_4696_p1);

assign add_ln700_220_fu_10456_p2 = (zext_ln142_344_fu_8433_p1 + zext_ln142_345_fu_8452_p1);

assign add_ln700_221_fu_10466_p2 = (zext_ln142_346_fu_8471_p1 + zext_ln142_347_fu_8490_p1);

assign add_ln700_222_fu_10476_p2 = (zext_ln700_216_fu_10472_p1 + zext_ln700_215_fu_10462_p1);

assign add_ln700_223_fu_10482_p2 = (zext_ln142_348_fu_8509_p1 + zext_ln142_349_fu_8528_p1);

assign add_ln700_224_fu_10492_p2 = (zext_ln142_350_fu_8547_p1 + zext_ln142_351_fu_8566_p1);

assign add_ln700_225_fu_10502_p2 = (zext_ln700_219_fu_10498_p1 + zext_ln700_218_fu_10488_p1);

assign add_ln700_226_fu_11358_p2 = (zext_ln700_220_fu_11355_p1 + zext_ln700_217_fu_11352_p1);

assign add_ln700_227_fu_10508_p2 = (zext_ln142_352_fu_8585_p1 + zext_ln142_353_fu_8604_p1);

assign add_ln700_228_fu_10518_p2 = (zext_ln142_354_fu_8623_p1 + zext_ln142_355_fu_8642_p1);

assign add_ln700_229_fu_10528_p2 = (zext_ln700_223_fu_10524_p1 + zext_ln700_222_fu_10514_p1);

assign add_ln700_22_fu_9166_p2 = (zext_ln142_48_fu_4719_p1 + zext_ln142_50_fu_4742_p1);

assign add_ln700_230_fu_10534_p2 = (zext_ln142_356_fu_8661_p1 + zext_ln142_357_fu_8680_p1);

assign add_ln700_231_fu_10544_p2 = (zext_ln142_358_fu_8699_p1 + zext_ln142_359_fu_8718_p1);

assign add_ln700_232_fu_10554_p2 = (zext_ln700_226_fu_10550_p1 + zext_ln700_225_fu_10540_p1);

assign add_ln700_233_fu_11374_p2 = (zext_ln700_227_fu_11371_p1 + zext_ln700_224_fu_11368_p1);

assign add_ln700_234_fu_11384_p2 = (zext_ln700_228_fu_11380_p1 + zext_ln700_221_fu_11364_p1);

assign add_ln700_235_fu_10560_p2 = (zext_ln142_360_fu_8737_p1 + zext_ln142_361_fu_8756_p1);

assign add_ln700_236_fu_10570_p2 = (zext_ln142_362_fu_8775_p1 + zext_ln142_363_fu_8794_p1);

assign add_ln700_237_fu_10580_p2 = (zext_ln700_231_fu_10576_p1 + zext_ln700_230_fu_10566_p1);

assign add_ln700_238_fu_10586_p2 = (zext_ln142_364_fu_8813_p1 + zext_ln142_365_fu_8832_p1);

assign add_ln700_239_fu_10596_p2 = (zext_ln142_366_fu_8851_p1 + zext_ln142_367_fu_8870_p1);

assign add_ln700_23_fu_9176_p2 = (zext_ln700_20_fu_9172_p1 + zext_ln700_19_fu_9162_p1);

assign add_ln700_240_fu_10606_p2 = (zext_ln700_234_fu_10602_p1 + zext_ln700_233_fu_10592_p1);

assign add_ln700_241_fu_11400_p2 = (zext_ln700_235_fu_11397_p1 + zext_ln700_232_fu_11394_p1);

assign add_ln700_242_fu_10612_p2 = (zext_ln142_368_fu_8889_p1 + zext_ln142_369_fu_8908_p1);

assign add_ln700_243_fu_10622_p2 = (zext_ln142_370_fu_8927_p1 + zext_ln142_371_fu_8946_p1);

assign add_ln700_244_fu_10632_p2 = (zext_ln700_238_fu_10628_p1 + zext_ln700_237_fu_10618_p1);

assign add_ln700_245_fu_10638_p2 = (zext_ln142_372_fu_8965_p1 + zext_ln142_373_fu_8984_p1);

assign add_ln700_246_fu_10648_p2 = (zext_ln142_374_fu_9003_p1 + zext_ln700_fu_9022_p1);

assign add_ln700_247_fu_10658_p2 = (zext_ln700_241_fu_10654_p1 + zext_ln700_240_fu_10644_p1);

assign add_ln700_248_fu_11416_p2 = (zext_ln700_242_fu_11413_p1 + zext_ln700_239_fu_11410_p1);

assign add_ln700_249_fu_11426_p2 = (zext_ln700_243_fu_11422_p1 + zext_ln700_236_fu_11406_p1);

assign add_ln700_24_fu_9182_p2 = (zext_ln142_52_fu_4765_p1 + zext_ln142_54_fu_4788_p1);

assign add_ln700_250_fu_11436_p2 = (zext_ln700_244_fu_11432_p1 + zext_ln700_229_fu_11390_p1);

assign add_ln700_251_fu_11446_p2 = (zext_ln700_245_fu_11442_p1 + zext_ln700_214_fu_11348_p1);

assign add_ln700_252_fu_11484_p2 = (zext_ln700_246_fu_11481_p1 + zext_ln700_183_fu_11478_p1);

assign add_ln700_25_fu_9192_p2 = (zext_ln142_56_fu_4811_p1 + zext_ln142_57_fu_4834_p1);

assign add_ln700_26_fu_9202_p2 = (zext_ln700_23_fu_9198_p1 + zext_ln700_22_fu_9188_p1);

assign add_ln700_27_fu_10764_p2 = (zext_ln700_24_fu_10761_p1 + zext_ln700_21_fu_10758_p1);

assign add_ln700_28_fu_10774_p2 = (zext_ln700_25_fu_10770_p1 + zext_ln700_18_fu_10754_p1);

assign add_ln700_29_fu_11455_p2 = (zext_ln700_26_fu_11452_p1 + add_ln700_13_reg_13375);

assign add_ln700_2_fu_9026_p2 = (zext_ln142_6_fu_4265_p1 + zext_ln142_8_fu_4284_p1);

assign add_ln700_30_fu_9208_p2 = (zext_ln142_59_fu_4853_p1 + zext_ln142_61_fu_4872_p1);

assign add_ln700_31_fu_9218_p2 = (zext_ln142_63_fu_4891_p1 + zext_ln142_65_fu_4910_p1);

assign add_ln700_32_fu_9228_p2 = (zext_ln700_28_fu_9224_p1 + zext_ln700_27_fu_9214_p1);

assign add_ln700_33_fu_9234_p2 = (zext_ln142_67_fu_4929_p1 + zext_ln142_69_fu_4948_p1);

assign add_ln700_34_fu_9244_p2 = (zext_ln142_71_fu_4967_p1 + zext_ln142_73_fu_4986_p1);

assign add_ln700_35_fu_9254_p2 = (zext_ln700_31_fu_9250_p1 + zext_ln700_30_fu_9240_p1);

assign add_ln700_36_fu_10786_p2 = (zext_ln700_32_fu_10783_p1 + zext_ln700_29_fu_10780_p1);

assign add_ln700_37_fu_9260_p2 = (zext_ln142_75_fu_5005_p1 + zext_ln142_77_fu_5024_p1);

assign add_ln700_38_fu_9270_p2 = (zext_ln142_79_fu_5043_p1 + zext_ln142_81_fu_5062_p1);

assign add_ln700_39_fu_9280_p2 = (zext_ln700_35_fu_9276_p1 + zext_ln700_34_fu_9266_p1);

assign add_ln700_3_fu_9036_p2 = (zext_ln142_10_fu_4307_p1 + zext_ln142_11_fu_4330_p1);

assign add_ln700_40_fu_9286_p2 = (zext_ln142_83_fu_5081_p1 + zext_ln142_85_fu_5100_p1);

assign add_ln700_41_fu_9296_p2 = (zext_ln142_87_fu_5119_p1 + zext_ln142_89_fu_5138_p1);

assign add_ln700_42_fu_9306_p2 = (zext_ln700_38_fu_9302_p1 + zext_ln700_37_fu_9292_p1);

assign add_ln700_43_fu_10802_p2 = (zext_ln700_39_fu_10799_p1 + zext_ln700_36_fu_10796_p1);

assign add_ln700_44_fu_10812_p2 = (zext_ln700_40_fu_10808_p1 + zext_ln700_33_fu_10792_p1);

assign add_ln700_45_fu_9312_p2 = (zext_ln142_91_fu_5161_p1 + zext_ln142_93_fu_5184_p1);

assign add_ln700_46_fu_9322_p2 = (zext_ln142_95_fu_5207_p1 + zext_ln142_97_fu_5230_p1);

assign add_ln700_47_fu_9332_p2 = (zext_ln700_43_fu_9328_p1 + zext_ln700_42_fu_9318_p1);

assign add_ln700_48_fu_9338_p2 = (zext_ln142_99_fu_5253_p1 + zext_ln142_101_fu_5276_p1);

assign add_ln700_49_fu_9348_p2 = (zext_ln142_103_fu_5299_p1 + zext_ln142_105_fu_5322_p1);

assign add_ln700_4_fu_9046_p2 = (zext_ln700_3_fu_9042_p1 + zext_ln700_2_fu_9032_p1);

assign add_ln700_50_fu_9358_p2 = (zext_ln700_46_fu_9354_p1 + zext_ln700_45_fu_9344_p1);

assign add_ln700_51_fu_10828_p2 = (zext_ln700_47_fu_10825_p1 + zext_ln700_44_fu_10822_p1);

assign add_ln700_52_fu_9364_p2 = (zext_ln142_107_fu_5345_p1 + zext_ln142_109_fu_5368_p1);

assign add_ln700_53_fu_9374_p2 = (zext_ln142_111_fu_5391_p1 + zext_ln142_113_fu_5414_p1);

assign add_ln700_54_fu_9384_p2 = (zext_ln700_50_fu_9380_p1 + zext_ln700_49_fu_9370_p1);

assign add_ln700_55_fu_9390_p2 = (zext_ln142_115_fu_5437_p1 + zext_ln142_117_fu_5460_p1);

assign add_ln700_56_fu_9400_p2 = (zext_ln142_119_fu_5483_p1 + zext_ln142_120_fu_5506_p1);

assign add_ln700_57_fu_9410_p2 = (zext_ln700_53_fu_9406_p1 + zext_ln700_52_fu_9396_p1);

assign add_ln700_58_fu_10844_p2 = (zext_ln700_54_fu_10841_p1 + zext_ln700_51_fu_10838_p1);

assign add_ln700_59_fu_10854_p2 = (zext_ln700_55_fu_10850_p1 + zext_ln700_48_fu_10834_p1);

assign add_ln700_5_fu_10714_p2 = (zext_ln700_4_fu_10711_p1 + add_ln700_1_fu_10705_p2);

assign add_ln700_60_fu_10864_p2 = (zext_ln700_56_fu_10860_p1 + zext_ln700_41_fu_10818_p1);

assign add_ln700_61_fu_11463_p2 = (zext_ln700_57_fu_11460_p1 + add_ln700_29_fu_11455_p2);

assign add_ln700_62_fu_9416_p2 = (zext_ln142_122_fu_5525_p1 + zext_ln142_124_fu_5544_p1);

assign add_ln700_63_fu_9426_p2 = (zext_ln142_126_fu_5563_p1 + zext_ln142_128_fu_5582_p1);

assign add_ln700_64_fu_9436_p2 = (zext_ln700_59_fu_9432_p1 + zext_ln700_58_fu_9422_p1);

assign add_ln700_65_fu_9442_p2 = (zext_ln142_130_fu_5601_p1 + zext_ln142_132_fu_5620_p1);

assign add_ln700_66_fu_9452_p2 = (zext_ln142_134_fu_5639_p1 + zext_ln142_136_fu_5658_p1);

assign add_ln700_67_fu_9462_p2 = (zext_ln700_62_fu_9458_p1 + zext_ln700_61_fu_9448_p1);

assign add_ln700_68_fu_10876_p2 = (zext_ln700_63_fu_10873_p1 + zext_ln700_60_fu_10870_p1);

assign add_ln700_69_fu_9468_p2 = (zext_ln142_138_fu_5677_p1 + zext_ln142_140_fu_5696_p1);

assign add_ln700_6_fu_9052_p2 = (zext_ln142_13_fu_4349_p1 + zext_ln142_15_fu_4368_p1);

assign add_ln700_70_fu_9478_p2 = (zext_ln142_142_fu_5715_p1 + zext_ln142_144_fu_5734_p1);

assign add_ln700_71_fu_9488_p2 = (zext_ln700_66_fu_9484_p1 + zext_ln700_65_fu_9474_p1);

assign add_ln700_72_fu_9494_p2 = (zext_ln142_146_fu_5753_p1 + zext_ln142_148_fu_5772_p1);

assign add_ln700_73_fu_9504_p2 = (zext_ln142_150_fu_5791_p1 + zext_ln142_152_fu_5810_p1);

assign add_ln700_74_fu_9514_p2 = (zext_ln700_69_fu_9510_p1 + zext_ln700_68_fu_9500_p1);

assign add_ln700_75_fu_10892_p2 = (zext_ln700_70_fu_10889_p1 + zext_ln700_67_fu_10886_p1);

assign add_ln700_76_fu_10902_p2 = (zext_ln700_71_fu_10898_p1 + zext_ln700_64_fu_10882_p1);

assign add_ln700_77_fu_9520_p2 = (zext_ln142_154_fu_5829_p1 + zext_ln142_156_fu_5848_p1);

assign add_ln700_78_fu_9530_p2 = (zext_ln142_158_fu_5867_p1 + zext_ln142_160_fu_5886_p1);

assign add_ln700_79_fu_9540_p2 = (zext_ln700_74_fu_9536_p1 + zext_ln700_73_fu_9526_p1);

assign add_ln700_7_fu_9062_p2 = (zext_ln142_17_fu_4387_p1 + zext_ln142_19_fu_4406_p1);

assign add_ln700_80_fu_9546_p2 = (zext_ln142_162_fu_5905_p1 + zext_ln142_164_fu_5924_p1);

assign add_ln700_81_fu_9556_p2 = (zext_ln142_166_fu_5943_p1 + zext_ln142_168_fu_5962_p1);

assign add_ln700_82_fu_9566_p2 = (zext_ln700_77_fu_9562_p1 + zext_ln700_76_fu_9552_p1);

assign add_ln700_83_fu_10918_p2 = (zext_ln700_78_fu_10915_p1 + zext_ln700_75_fu_10912_p1);

assign add_ln700_84_fu_9572_p2 = (zext_ln142_170_fu_5981_p1 + zext_ln142_172_fu_6000_p1);

assign add_ln700_85_fu_9582_p2 = (zext_ln142_174_fu_6019_p1 + zext_ln142_176_fu_6038_p1);

assign add_ln700_86_fu_9592_p2 = (zext_ln700_81_fu_9588_p1 + zext_ln700_80_fu_9578_p1);

assign add_ln700_87_fu_9598_p2 = (zext_ln142_178_fu_6057_p1 + zext_ln142_180_fu_6076_p1);

assign add_ln700_88_fu_9608_p2 = (zext_ln142_182_fu_6095_p1 + zext_ln142_184_fu_6114_p1);

assign add_ln700_89_fu_9618_p2 = (zext_ln700_84_fu_9614_p1 + zext_ln700_83_fu_9604_p1);

assign add_ln700_8_fu_9072_p2 = (zext_ln700_6_fu_9068_p1 + zext_ln700_5_fu_9058_p1);

assign add_ln700_90_fu_10934_p2 = (zext_ln700_85_fu_10931_p1 + zext_ln700_82_fu_10928_p1);

assign add_ln700_91_fu_10944_p2 = (zext_ln700_86_fu_10940_p1 + zext_ln700_79_fu_10924_p1);

assign add_ln700_92_fu_10954_p2 = (zext_ln700_87_fu_10950_p1 + zext_ln700_72_fu_10908_p1);

assign add_ln700_93_fu_9624_p2 = (zext_ln142_186_fu_6137_p1 + zext_ln142_188_fu_6160_p1);

assign add_ln700_94_fu_9634_p2 = (zext_ln142_190_fu_6183_p1 + zext_ln142_192_fu_6206_p1);

assign add_ln700_95_fu_9644_p2 = (zext_ln700_90_fu_9640_p1 + zext_ln700_89_fu_9630_p1);

assign add_ln700_96_fu_9650_p2 = (zext_ln142_194_fu_6229_p1 + zext_ln142_196_fu_6252_p1);

assign add_ln700_97_fu_9660_p2 = (zext_ln142_198_fu_6275_p1 + zext_ln142_200_fu_6298_p1);

assign add_ln700_98_fu_9670_p2 = (zext_ln700_93_fu_9666_p1 + zext_ln700_92_fu_9656_p1);

assign add_ln700_99_fu_10970_p2 = (zext_ln700_94_fu_10967_p1 + zext_ln700_91_fu_10964_p1);

assign add_ln700_9_fu_9078_p2 = (zext_ln142_21_fu_4429_p1 + zext_ln142_23_fu_4452_p1);

assign add_ln700_fu_10695_p2 = (zext_ln142_3_fu_10682_p1 + zext_ln142_4_fu_10691_p1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state6 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_3928_p2 == 1'd0));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_block_state5_io)) | ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_3928_p2 == 1'd0)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_block_state5_io)) | ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_3928_p2 == 1'd0)));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = ((in_V_V_TVALID == 1'b0) & (icmp_ln221_fu_3928_p2 == 1'd0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state5_io = ((out_V_V_TREADY == 1'b0) & (icmp_ln221_reg_11497_pp0_iter2_reg == 1'd0));
end

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign i_fu_3934_p2 = (i_0_reg_3917 + 12'd1);

assign icmp_ln221_fu_3928_p2 = ((i_0_reg_3917 == 12'd3072) ? 1'b1 : 1'b0);

assign icmp_ln235_fu_4205_p2 = ((nf_fu_4199_p2 == 32'd3) ? 1'b1 : 1'b0);

assign icmp_ln899_100_fu_6241_p2 = ((tmp_V_1_reg_11506 < zext_ln142_195_fu_6237_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_101_fu_6264_p2 = ((tmp_V_1_reg_11506 < zext_ln142_197_fu_6260_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_102_fu_6287_p2 = ((tmp_V_1_reg_11506 < zext_ln142_199_fu_6283_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_103_fu_6310_p2 = ((tmp_V_1_reg_11506 < zext_ln142_201_fu_6306_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_104_fu_6333_p2 = ((tmp_V_1_reg_11506 < zext_ln142_203_fu_6329_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_105_fu_6356_p2 = ((tmp_V_1_reg_11506 < zext_ln142_205_fu_6352_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_106_fu_6379_p2 = ((tmp_V_1_reg_11506 < zext_ln142_207_fu_6375_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_107_fu_6402_p2 = ((tmp_V_1_reg_11506 < zext_ln142_209_fu_6398_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_108_fu_6425_p2 = ((tmp_V_1_reg_11506 < zext_ln142_211_fu_6421_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_109_fu_6448_p2 = ((tmp_V_1_reg_11506 < zext_ln142_213_fu_6444_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_10_fu_4395_p2 = ((tmp_V_1_reg_11506 < zext_ln142_18_fu_4391_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_110_fu_6471_p2 = ((tmp_V_1_reg_11506 < zext_ln142_215_fu_6467_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_111_fu_6494_p2 = ((tmp_V_1_reg_11506 < zext_ln142_217_fu_6490_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_112_fu_6517_p2 = ((tmp_V_1_reg_11506 < zext_ln142_219_fu_6513_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_113_fu_6540_p2 = ((tmp_V_1_reg_11506 < zext_ln142_221_fu_6536_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_114_fu_6563_p2 = ((tmp_V_1_reg_11506 < zext_ln142_223_fu_6559_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_115_fu_6586_p2 = ((tmp_V_1_reg_11506 < zext_ln142_225_fu_6582_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_116_fu_6609_p2 = ((tmp_V_1_reg_11506 < zext_ln142_227_fu_6605_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_117_fu_6632_p2 = ((tmp_V_1_reg_11506 < zext_ln142_229_fu_6628_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_118_fu_6655_p2 = ((tmp_V_1_reg_11506 < zext_ln142_231_fu_6651_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_119_fu_6678_p2 = ((tmp_V_1_reg_11506 < zext_ln142_233_fu_6674_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_11_fu_4418_p2 = ((tmp_V_1_reg_11506 < zext_ln142_20_fu_4414_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_120_fu_6701_p2 = ((tmp_V_1_reg_11506 < zext_ln142_235_fu_6697_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_121_fu_6724_p2 = ((tmp_V_1_reg_11506 < zext_ln142_237_fu_6720_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_122_fu_6747_p2 = ((tmp_V_1_reg_11506 < zext_ln142_239_fu_6743_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_123_fu_6770_p2 = ((tmp_V_1_reg_11506 < zext_ln142_241_fu_6766_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_124_fu_6793_p2 = ((tmp_V_1_reg_11506 < zext_ln142_243_fu_6789_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_125_fu_6816_p2 = ((tmp_V_1_reg_11506 < zext_ln142_245_fu_6812_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_126_fu_6839_p2 = ((tmp_V_1_reg_11506 < select_ln142_5_fu_6831_p3) ? 1'b1 : 1'b0);

assign icmp_ln899_127_fu_6854_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_222_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_128_fu_6869_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_221_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_129_fu_6884_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_220_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_12_fu_4441_p2 = ((tmp_V_1_reg_11506 < zext_ln142_22_fu_4437_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_130_fu_6899_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_218_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_131_fu_6914_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_217_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_132_fu_6929_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_216_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_133_fu_6944_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_215_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_134_fu_6959_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_214_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_135_fu_6974_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_213_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_136_fu_6989_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_212_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_137_fu_7004_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_211_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_138_fu_7019_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_210_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_139_fu_7034_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_209_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_13_fu_4464_p2 = ((tmp_V_1_reg_11506 < zext_ln142_24_fu_4460_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_140_fu_7049_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_207_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_141_fu_7064_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_206_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_142_fu_7079_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_205_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_143_fu_7094_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_204_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_144_fu_7109_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_203_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_145_fu_7124_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_202_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_146_fu_7139_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_201_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_147_fu_7154_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_200_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_148_fu_7169_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_199_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_149_fu_7184_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_198_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_14_fu_4487_p2 = ((tmp_V_1_reg_11506 < select_ln142_2_fu_4479_p3) ? 1'b1 : 1'b0);

assign icmp_ln899_150_fu_7199_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_196_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_151_fu_7214_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_195_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_152_fu_7229_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_194_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_153_fu_7244_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_193_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_154_fu_7259_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_192_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_155_fu_7274_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_191_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_156_fu_7289_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_190_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_157_fu_7304_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_189_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_158_fu_7319_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_188_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_159_fu_7334_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_187_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_15_fu_4506_p2 = ((tmp_V_1_reg_11506 < zext_ln142_27_fu_4502_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_160_fu_7349_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_185_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_161_fu_7364_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_184_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_162_fu_7379_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_183_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_163_fu_7394_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_182_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_164_fu_7409_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_181_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_165_fu_7424_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_180_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_166_fu_7439_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_179_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_167_fu_7454_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_178_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_168_fu_7469_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_177_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_169_fu_7484_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_176_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_16_fu_4525_p2 = ((tmp_V_1_reg_11506 < zext_ln142_29_fu_4521_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_170_fu_7499_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_174_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_171_fu_7514_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_173_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_172_fu_7529_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_172_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_173_fu_7544_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_171_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_174_fu_7559_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_170_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_175_fu_7574_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_169_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_176_fu_7589_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_168_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_177_fu_7604_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_167_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_178_fu_7619_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_166_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_179_fu_7634_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_165_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_17_fu_4544_p2 = ((tmp_V_1_reg_11506 < zext_ln142_31_fu_4540_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_180_fu_7649_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_163_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_181_fu_7664_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_162_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_182_fu_7679_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_161_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_183_fu_7694_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_160_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_184_fu_7709_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_159_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_185_fu_7724_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_158_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_186_fu_7739_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_157_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_187_fu_7754_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_156_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_188_fu_7769_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_155_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_189_fu_7784_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_154_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_18_fu_4563_p2 = ((tmp_V_1_reg_11506 < zext_ln142_33_fu_4559_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_190_fu_7799_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_152_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_191_fu_7814_p2 = ((tmp_V_1_reg_11506 < threshs_m_thresholds_151_q0) ? 1'b1 : 1'b0);

assign icmp_ln899_192_fu_7833_p2 = ((tmp_V_1_reg_11506 < sext_ln142_57_fu_7829_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_193_fu_7852_p2 = ((tmp_V_1_reg_11506 < sext_ln142_58_fu_7848_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_194_fu_7871_p2 = ((tmp_V_1_reg_11506 < sext_ln142_59_fu_7867_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_195_fu_7890_p2 = ((tmp_V_1_reg_11506 < sext_ln142_60_fu_7886_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_196_fu_7909_p2 = ((tmp_V_1_reg_11506 < sext_ln142_61_fu_7905_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_197_fu_7928_p2 = ((tmp_V_1_reg_11506 < sext_ln142_62_fu_7924_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_198_fu_7947_p2 = ((tmp_V_1_reg_11506 < sext_ln142_63_fu_7943_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_199_fu_7966_p2 = ((tmp_V_1_reg_11506 < sext_ln142_64_fu_7962_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_19_fu_4582_p2 = ((tmp_V_1_reg_11506 < zext_ln142_35_fu_4578_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_1_fu_4232_p2 = ((tmp_V_1_reg_11506 < zext_ln142_2_fu_4228_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_200_fu_7985_p2 = ((tmp_V_1_reg_11506 < sext_ln142_65_fu_7981_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_201_fu_8004_p2 = ((tmp_V_1_reg_11506 < sext_ln142_66_fu_8000_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_202_fu_8023_p2 = ((tmp_V_1_reg_11506 < sext_ln142_67_fu_8019_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_203_fu_8042_p2 = ((tmp_V_1_reg_11506 < sext_ln142_68_fu_8038_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_204_fu_8061_p2 = ((tmp_V_1_reg_11506 < sext_ln142_69_fu_8057_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_205_fu_8080_p2 = ((tmp_V_1_reg_11506 < sext_ln142_70_fu_8076_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_206_fu_8099_p2 = ((tmp_V_1_reg_11506 < sext_ln142_71_fu_8095_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_207_fu_8118_p2 = ((tmp_V_1_reg_11506 < sext_ln142_72_fu_8114_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_208_fu_8137_p2 = ((tmp_V_1_reg_11506 < sext_ln142_73_fu_8133_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_209_fu_8156_p2 = ((tmp_V_1_reg_11506 < sext_ln142_74_fu_8152_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_20_fu_4601_p2 = ((tmp_V_1_reg_11506 < zext_ln142_37_fu_4597_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_210_fu_8175_p2 = ((tmp_V_1_reg_11506 < sext_ln142_75_fu_8171_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_211_fu_8194_p2 = ((tmp_V_1_reg_11506 < sext_ln142_76_fu_8190_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_212_fu_8213_p2 = ((tmp_V_1_reg_11506 < sext_ln142_77_fu_8209_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_213_fu_8232_p2 = ((tmp_V_1_reg_11506 < sext_ln142_78_fu_8228_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_214_fu_8251_p2 = ((tmp_V_1_reg_11506 < sext_ln142_79_fu_8247_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_215_fu_8270_p2 = ((tmp_V_1_reg_11506 < sext_ln142_80_fu_8266_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_216_fu_8289_p2 = ((tmp_V_1_reg_11506 < sext_ln142_81_fu_8285_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_217_fu_8308_p2 = ((tmp_V_1_reg_11506 < sext_ln142_82_fu_8304_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_218_fu_8327_p2 = ((tmp_V_1_reg_11506 < sext_ln142_83_fu_8323_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_219_fu_8346_p2 = ((tmp_V_1_reg_11506 < sext_ln142_84_fu_8342_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_21_fu_4620_p2 = ((tmp_V_1_reg_11506 < zext_ln142_39_fu_4616_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_220_fu_8365_p2 = ((tmp_V_1_reg_11506 < sext_ln142_85_fu_8361_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_221_fu_8384_p2 = ((tmp_V_1_reg_11506 < sext_ln142_86_fu_8380_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_222_fu_8403_p2 = ((tmp_V_1_reg_11506 < sext_ln142_87_fu_8399_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_223_fu_8422_p2 = ((tmp_V_1_reg_11506 < sext_ln142_88_fu_8418_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_224_fu_8441_p2 = ((tmp_V_1_reg_11506 < sext_ln142_89_fu_8437_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_225_fu_8460_p2 = ((tmp_V_1_reg_11506 < sext_ln142_90_fu_8456_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_226_fu_8479_p2 = ((tmp_V_1_reg_11506 < sext_ln142_91_fu_8475_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_227_fu_8498_p2 = ((tmp_V_1_reg_11506 < sext_ln142_92_fu_8494_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_228_fu_8517_p2 = ((tmp_V_1_reg_11506 < sext_ln142_93_fu_8513_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_229_fu_8536_p2 = ((tmp_V_1_reg_11506 < sext_ln142_94_fu_8532_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_22_fu_4639_p2 = ((tmp_V_1_reg_11506 < zext_ln142_41_fu_4635_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_230_fu_8555_p2 = ((tmp_V_1_reg_11506 < sext_ln142_95_fu_8551_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_231_fu_8574_p2 = ((tmp_V_1_reg_11506 < sext_ln142_96_fu_8570_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_232_fu_8593_p2 = ((tmp_V_1_reg_11506 < sext_ln142_97_fu_8589_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_233_fu_8612_p2 = ((tmp_V_1_reg_11506 < sext_ln142_98_fu_8608_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_234_fu_8631_p2 = ((tmp_V_1_reg_11506 < sext_ln142_99_fu_8627_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_235_fu_8650_p2 = ((tmp_V_1_reg_11506 < sext_ln142_100_fu_8646_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_236_fu_8669_p2 = ((tmp_V_1_reg_11506 < sext_ln142_101_fu_8665_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_237_fu_8688_p2 = ((tmp_V_1_reg_11506 < sext_ln142_102_fu_8684_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_238_fu_8707_p2 = ((tmp_V_1_reg_11506 < sext_ln142_103_fu_8703_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_239_fu_8726_p2 = ((tmp_V_1_reg_11506 < sext_ln142_104_fu_8722_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_23_fu_4662_p2 = ((tmp_V_1_reg_11506 < zext_ln142_43_fu_4658_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_240_fu_8745_p2 = ((tmp_V_1_reg_11506 < sext_ln142_105_fu_8741_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_241_fu_8764_p2 = ((tmp_V_1_reg_11506 < sext_ln142_106_fu_8760_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_242_fu_8783_p2 = ((tmp_V_1_reg_11506 < sext_ln142_107_fu_8779_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_243_fu_8802_p2 = ((tmp_V_1_reg_11506 < sext_ln142_108_fu_8798_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_244_fu_8821_p2 = ((tmp_V_1_reg_11506 < sext_ln142_109_fu_8817_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_245_fu_8840_p2 = ((tmp_V_1_reg_11506 < sext_ln142_110_fu_8836_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_246_fu_8859_p2 = ((tmp_V_1_reg_11506 < sext_ln142_111_fu_8855_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_247_fu_8878_p2 = ((tmp_V_1_reg_11506 < sext_ln142_112_fu_8874_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_248_fu_8897_p2 = ((tmp_V_1_reg_11506 < sext_ln142_113_fu_8893_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_249_fu_8916_p2 = ((tmp_V_1_reg_11506 < sext_ln142_114_fu_8912_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_24_fu_4685_p2 = ((tmp_V_1_reg_11506 < zext_ln142_45_fu_4681_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_250_fu_8935_p2 = ((tmp_V_1_reg_11506 < sext_ln142_115_fu_8931_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_251_fu_8954_p2 = ((tmp_V_1_reg_11506 < sext_ln142_116_fu_8950_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_252_fu_8973_p2 = ((tmp_V_1_reg_11506 < sext_ln142_117_fu_8969_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_253_fu_8992_p2 = ((tmp_V_1_reg_11506 < sext_ln142_118_fu_8988_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_254_fu_9011_p2 = ((tmp_V_1_reg_11506 < sext_ln142_119_fu_9007_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_25_fu_4708_p2 = ((tmp_V_1_reg_11506 < zext_ln142_47_fu_4704_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_26_fu_4731_p2 = ((tmp_V_1_reg_11506 < zext_ln142_49_fu_4727_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_27_fu_4754_p2 = ((tmp_V_1_reg_11506 < zext_ln142_51_fu_4750_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_28_fu_4777_p2 = ((tmp_V_1_reg_11506 < zext_ln142_53_fu_4773_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_29_fu_4800_p2 = ((tmp_V_1_reg_11506 < zext_ln142_55_fu_4796_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_2_fu_4245_p2 = ((tmp_V_1_reg_11506 < select_ln142_fu_4237_p3) ? 1'b1 : 1'b0);

assign icmp_ln899_30_fu_4823_p2 = ((tmp_V_1_reg_11506 < select_ln142_3_fu_4815_p3) ? 1'b1 : 1'b0);

assign icmp_ln899_31_fu_4842_p2 = ((tmp_V_1_reg_11506 < zext_ln142_58_fu_4838_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_32_fu_4861_p2 = ((tmp_V_1_reg_11506 < zext_ln142_60_fu_4857_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_33_fu_4880_p2 = ((tmp_V_1_reg_11506 < zext_ln142_62_fu_4876_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_34_fu_4899_p2 = ((tmp_V_1_reg_11506 < zext_ln142_64_fu_4895_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_35_fu_4918_p2 = ((tmp_V_1_reg_11506 < zext_ln142_66_fu_4914_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_36_fu_4937_p2 = ((tmp_V_1_reg_11506 < zext_ln142_68_fu_4933_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_37_fu_4956_p2 = ((tmp_V_1_reg_11506 < zext_ln142_70_fu_4952_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_38_fu_4975_p2 = ((tmp_V_1_reg_11506 < zext_ln142_72_fu_4971_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_39_fu_4994_p2 = ((tmp_V_1_reg_11506 < zext_ln142_74_fu_4990_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_3_fu_4254_p2 = ((tmp_V_1_reg_11506 < zext_ln142_5_fu_4250_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_40_fu_5013_p2 = ((tmp_V_1_reg_11506 < zext_ln142_76_fu_5009_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_41_fu_5032_p2 = ((tmp_V_1_reg_11506 < zext_ln142_78_fu_5028_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_42_fu_5051_p2 = ((tmp_V_1_reg_11506 < zext_ln142_80_fu_5047_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_43_fu_5070_p2 = ((tmp_V_1_reg_11506 < zext_ln142_82_fu_5066_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_44_fu_5089_p2 = ((tmp_V_1_reg_11506 < zext_ln142_84_fu_5085_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_45_fu_5108_p2 = ((tmp_V_1_reg_11506 < zext_ln142_86_fu_5104_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_46_fu_5127_p2 = ((tmp_V_1_reg_11506 < zext_ln142_88_fu_5123_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_47_fu_5150_p2 = ((tmp_V_1_reg_11506 < zext_ln142_90_fu_5146_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_48_fu_5173_p2 = ((tmp_V_1_reg_11506 < zext_ln142_92_fu_5169_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_49_fu_5196_p2 = ((tmp_V_1_reg_11506 < zext_ln142_94_fu_5192_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_4_fu_4273_p2 = ((tmp_V_1_reg_11506 < zext_ln142_7_fu_4269_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_50_fu_5219_p2 = ((tmp_V_1_reg_11506 < zext_ln142_96_fu_5215_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_51_fu_5242_p2 = ((tmp_V_1_reg_11506 < zext_ln142_98_fu_5238_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_52_fu_5265_p2 = ((tmp_V_1_reg_11506 < zext_ln142_100_fu_5261_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_53_fu_5288_p2 = ((tmp_V_1_reg_11506 < zext_ln142_102_fu_5284_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_54_fu_5311_p2 = ((tmp_V_1_reg_11506 < zext_ln142_104_fu_5307_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_55_fu_5334_p2 = ((tmp_V_1_reg_11506 < zext_ln142_106_fu_5330_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_56_fu_5357_p2 = ((tmp_V_1_reg_11506 < zext_ln142_108_fu_5353_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_57_fu_5380_p2 = ((tmp_V_1_reg_11506 < zext_ln142_110_fu_5376_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_58_fu_5403_p2 = ((tmp_V_1_reg_11506 < zext_ln142_112_fu_5399_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_59_fu_5426_p2 = ((tmp_V_1_reg_11506 < zext_ln142_114_fu_5422_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_5_fu_4296_p2 = ((tmp_V_1_reg_11506 < zext_ln142_9_fu_4292_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_60_fu_5449_p2 = ((tmp_V_1_reg_11506 < zext_ln142_116_fu_5445_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_61_fu_5472_p2 = ((tmp_V_1_reg_11506 < zext_ln142_118_fu_5468_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_62_fu_5495_p2 = ((tmp_V_1_reg_11506 < select_ln142_4_fu_5487_p3) ? 1'b1 : 1'b0);

assign icmp_ln899_63_fu_5514_p2 = ((tmp_V_1_reg_11506 < zext_ln142_121_fu_5510_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_64_fu_5533_p2 = ((tmp_V_1_reg_11506 < zext_ln142_123_fu_5529_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_65_fu_5552_p2 = ((tmp_V_1_reg_11506 < zext_ln142_125_fu_5548_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_66_fu_5571_p2 = ((tmp_V_1_reg_11506 < zext_ln142_127_fu_5567_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_67_fu_5590_p2 = ((tmp_V_1_reg_11506 < zext_ln142_129_fu_5586_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_68_fu_5609_p2 = ((tmp_V_1_reg_11506 < zext_ln142_131_fu_5605_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_69_fu_5628_p2 = ((tmp_V_1_reg_11506 < zext_ln142_133_fu_5624_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_6_fu_4319_p2 = ((tmp_V_1_reg_11506 < select_ln142_1_fu_4311_p3) ? 1'b1 : 1'b0);

assign icmp_ln899_70_fu_5647_p2 = ((tmp_V_1_reg_11506 < zext_ln142_135_fu_5643_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_71_fu_5666_p2 = ((tmp_V_1_reg_11506 < zext_ln142_137_fu_5662_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_72_fu_5685_p2 = ((tmp_V_1_reg_11506 < zext_ln142_139_fu_5681_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_73_fu_5704_p2 = ((tmp_V_1_reg_11506 < zext_ln142_141_fu_5700_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_74_fu_5723_p2 = ((tmp_V_1_reg_11506 < zext_ln142_143_fu_5719_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_75_fu_5742_p2 = ((tmp_V_1_reg_11506 < zext_ln142_145_fu_5738_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_76_fu_5761_p2 = ((tmp_V_1_reg_11506 < zext_ln142_147_fu_5757_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_77_fu_5780_p2 = ((tmp_V_1_reg_11506 < zext_ln142_149_fu_5776_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_78_fu_5799_p2 = ((tmp_V_1_reg_11506 < zext_ln142_151_fu_5795_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_79_fu_5818_p2 = ((tmp_V_1_reg_11506 < zext_ln142_153_fu_5814_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_7_fu_4338_p2 = ((tmp_V_1_reg_11506 < zext_ln142_12_fu_4334_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_80_fu_5837_p2 = ((tmp_V_1_reg_11506 < zext_ln142_155_fu_5833_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_81_fu_5856_p2 = ((tmp_V_1_reg_11506 < zext_ln142_157_fu_5852_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_82_fu_5875_p2 = ((tmp_V_1_reg_11506 < zext_ln142_159_fu_5871_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_83_fu_5894_p2 = ((tmp_V_1_reg_11506 < zext_ln142_161_fu_5890_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_84_fu_5913_p2 = ((tmp_V_1_reg_11506 < zext_ln142_163_fu_5909_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_85_fu_5932_p2 = ((tmp_V_1_reg_11506 < zext_ln142_165_fu_5928_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_86_fu_5951_p2 = ((tmp_V_1_reg_11506 < zext_ln142_167_fu_5947_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_87_fu_5970_p2 = ((tmp_V_1_reg_11506 < zext_ln142_169_fu_5966_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_88_fu_5989_p2 = ((tmp_V_1_reg_11506 < zext_ln142_171_fu_5985_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_89_fu_6008_p2 = ((tmp_V_1_reg_11506 < zext_ln142_173_fu_6004_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_8_fu_4357_p2 = ((tmp_V_1_reg_11506 < zext_ln142_14_fu_4353_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_90_fu_6027_p2 = ((tmp_V_1_reg_11506 < zext_ln142_175_fu_6023_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_91_fu_6046_p2 = ((tmp_V_1_reg_11506 < zext_ln142_177_fu_6042_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_92_fu_6065_p2 = ((tmp_V_1_reg_11506 < zext_ln142_179_fu_6061_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_93_fu_6084_p2 = ((tmp_V_1_reg_11506 < zext_ln142_181_fu_6080_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_94_fu_6103_p2 = ((tmp_V_1_reg_11506 < zext_ln142_183_fu_6099_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_95_fu_6126_p2 = ((tmp_V_1_reg_11506 < zext_ln142_185_fu_6122_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_96_fu_6149_p2 = ((tmp_V_1_reg_11506 < zext_ln142_187_fu_6145_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_97_fu_6172_p2 = ((tmp_V_1_reg_11506 < zext_ln142_189_fu_6168_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_98_fu_6195_p2 = ((tmp_V_1_reg_11506 < zext_ln142_191_fu_6191_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_99_fu_6218_p2 = ((tmp_V_1_reg_11506 < zext_ln142_193_fu_6214_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_9_fu_4376_p2 = ((tmp_V_1_reg_11506 < zext_ln142_16_fu_4372_p1) ? 1'b1 : 1'b0);

assign icmp_ln899_fu_4223_p2 = ((tmp_V_1_reg_11506 < zext_ln142_1_fu_4219_p1) ? 1'b1 : 1'b0);

assign nf_1_fu_4211_p3 = ((icmp_ln235_fu_4205_p2[0:0] === 1'b1) ? 32'd0 : nf_fu_4199_p2);

assign nf_fu_4199_p2 = (nf_assign_reg_3906 + 32'd1);

assign or_ln_fu_10669_p3 = {{7'd64}, {xor_ln899_fu_10664_p2}};

assign out_V_V_TDATA = (add_ln700_252_fu_11484_p2 + add_ln700_125_fu_11472_p2);

assign select_ln142_1_fu_4311_p3 = ((threshs_m_thresholds_43_q0[0:0] === 1'b1) ? 8'd7 : 8'd0);

assign select_ln142_2_fu_4479_p3 = ((threshs_m_thresholds_208_q0[0:0] === 1'b1) ? 8'd15 : 8'd0);

assign select_ln142_3_fu_4815_p3 = ((threshs_m_thresholds_75_q0[0:0] === 1'b1) ? 8'd31 : 8'd0);

assign select_ln142_4_fu_5487_p3 = ((threshs_m_thresholds_40_q0[0:0] === 1'b1) ? 8'd63 : 8'd0);

assign select_ln142_5_fu_6831_p3 = ((threshs_m_thresholds_223_q0[0:0] === 1'b1) ? 8'd127 : 8'd0);

assign select_ln142_fu_4237_p3 = ((threshs_m_thresholds_142_q0[0:0] === 1'b1) ? 8'd3 : 8'd0);

assign sext_ln142_100_fu_8646_p1 = $signed(threshs_m_thresholds_102_q0);

assign sext_ln142_101_fu_8665_p1 = $signed(threshs_m_thresholds_101_q0);

assign sext_ln142_102_fu_8684_p1 = $signed(threshs_m_thresholds_100_q0);

assign sext_ln142_103_fu_8703_p1 = $signed(threshs_m_thresholds_99_q0);

assign sext_ln142_104_fu_8722_p1 = $signed(threshs_m_thresholds_98_q0);

assign sext_ln142_105_fu_8741_p1 = $signed(threshs_m_thresholds_96_q0);

assign sext_ln142_106_fu_8760_p1 = $signed(threshs_m_thresholds_95_q0);

assign sext_ln142_107_fu_8779_p1 = $signed(threshs_m_thresholds_94_q0);

assign sext_ln142_108_fu_8798_p1 = $signed(threshs_m_thresholds_93_q0);

assign sext_ln142_109_fu_8817_p1 = $signed(threshs_m_thresholds_92_q0);

assign sext_ln142_10_fu_4792_p1 = $signed(threshs_m_thresholds_77_q0);

assign sext_ln142_110_fu_8836_p1 = $signed(threshs_m_thresholds_91_q0);

assign sext_ln142_111_fu_8855_p1 = $signed(threshs_m_thresholds_90_q0);

assign sext_ln142_112_fu_8874_p1 = $signed(threshs_m_thresholds_89_q0);

assign sext_ln142_113_fu_8893_p1 = $signed(threshs_m_thresholds_88_q0);

assign sext_ln142_114_fu_8912_p1 = $signed(threshs_m_thresholds_87_q0);

assign sext_ln142_115_fu_8931_p1 = $signed(threshs_m_thresholds_85_q0);

assign sext_ln142_116_fu_8950_p1 = $signed(threshs_m_thresholds_84_q0);

assign sext_ln142_117_fu_8969_p1 = $signed(threshs_m_thresholds_83_q0);

assign sext_ln142_118_fu_8988_p1 = $signed(threshs_m_thresholds_82_q0);

assign sext_ln142_119_fu_9007_p1 = $signed(threshs_m_thresholds_81_q0);

assign sext_ln142_11_fu_5142_p1 = $signed(threshs_m_thresholds_57_q0);

assign sext_ln142_12_fu_5165_p1 = $signed(threshs_m_thresholds_56_q0);

assign sext_ln142_13_fu_5188_p1 = $signed(threshs_m_thresholds_55_q0);

assign sext_ln142_14_fu_5211_p1 = $signed(threshs_m_thresholds_53_q0);

assign sext_ln142_15_fu_5234_p1 = $signed(threshs_m_thresholds_52_q0);

assign sext_ln142_16_fu_5257_p1 = $signed(threshs_m_thresholds_51_q0);

assign sext_ln142_17_fu_5280_p1 = $signed(threshs_m_thresholds_50_q0);

assign sext_ln142_18_fu_5303_p1 = $signed(threshs_m_thresholds_49_q0);

assign sext_ln142_19_fu_5326_p1 = $signed(threshs_m_thresholds_48_q0);

assign sext_ln142_1_fu_4410_p1 = $signed(threshs_m_thresholds_241_q0);

assign sext_ln142_20_fu_5349_p1 = $signed(threshs_m_thresholds_47_q0);

assign sext_ln142_21_fu_5372_p1 = $signed(threshs_m_thresholds_46_q0);

assign sext_ln142_22_fu_5395_p1 = $signed(threshs_m_thresholds_45_q0);

assign sext_ln142_23_fu_5418_p1 = $signed(threshs_m_thresholds_44_q0);

assign sext_ln142_24_fu_5441_p1 = $signed(threshs_m_thresholds_42_q0);

assign sext_ln142_25_fu_5464_p1 = $signed(threshs_m_thresholds_41_q0);

assign sext_ln142_26_fu_6118_p1 = $signed(threshs_m_thresholds_4_q0);

assign sext_ln142_27_fu_6141_p1 = $signed(threshs_m_thresholds_3_q0);

assign sext_ln142_28_fu_6164_p1 = $signed(threshs_m_thresholds_2_q0);

assign sext_ln142_29_fu_6187_p1 = $signed(threshs_m_thresholds_1_q0);

assign sext_ln142_2_fu_4433_p1 = $signed(threshs_m_thresholds_230_q0);

assign sext_ln142_30_fu_6210_p1 = $signed(threshs_m_thresholds_q0);

assign sext_ln142_31_fu_6233_p1 = $signed(threshs_m_thresholds_251_q0);

assign sext_ln142_32_fu_6256_p1 = $signed(threshs_m_thresholds_250_q0);

assign sext_ln142_33_fu_6279_p1 = $signed(threshs_m_thresholds_249_q0);

assign sext_ln142_34_fu_6302_p1 = $signed(threshs_m_thresholds_248_q0);

assign sext_ln142_35_fu_6325_p1 = $signed(threshs_m_thresholds_247_q0);

assign sext_ln142_36_fu_6348_p1 = $signed(threshs_m_thresholds_246_q0);

assign sext_ln142_37_fu_6371_p1 = $signed(threshs_m_thresholds_245_q0);

assign sext_ln142_38_fu_6394_p1 = $signed(threshs_m_thresholds_244_q0);

assign sext_ln142_39_fu_6417_p1 = $signed(threshs_m_thresholds_243_q0);

assign sext_ln142_3_fu_4456_p1 = $signed(threshs_m_thresholds_219_q0);

assign sext_ln142_40_fu_6440_p1 = $signed(threshs_m_thresholds_242_q0);

assign sext_ln142_41_fu_6463_p1 = $signed(threshs_m_thresholds_240_q0);

assign sext_ln142_42_fu_6486_p1 = $signed(threshs_m_thresholds_239_q0);

assign sext_ln142_43_fu_6509_p1 = $signed(threshs_m_thresholds_238_q0);

assign sext_ln142_44_fu_6532_p1 = $signed(threshs_m_thresholds_237_q0);

assign sext_ln142_45_fu_6555_p1 = $signed(threshs_m_thresholds_236_q0);

assign sext_ln142_46_fu_6578_p1 = $signed(threshs_m_thresholds_235_q0);

assign sext_ln142_47_fu_6601_p1 = $signed(threshs_m_thresholds_234_q0);

assign sext_ln142_48_fu_6624_p1 = $signed(threshs_m_thresholds_233_q0);

assign sext_ln142_49_fu_6647_p1 = $signed(threshs_m_thresholds_232_q0);

assign sext_ln142_4_fu_4654_p1 = $signed(threshs_m_thresholds_108_q0);

assign sext_ln142_50_fu_6670_p1 = $signed(threshs_m_thresholds_231_q0);

assign sext_ln142_51_fu_6693_p1 = $signed(threshs_m_thresholds_229_q0);

assign sext_ln142_52_fu_6716_p1 = $signed(threshs_m_thresholds_228_q0);

assign sext_ln142_53_fu_6739_p1 = $signed(threshs_m_thresholds_227_q0);

assign sext_ln142_54_fu_6762_p1 = $signed(threshs_m_thresholds_226_q0);

assign sext_ln142_55_fu_6785_p1 = $signed(threshs_m_thresholds_225_q0);

assign sext_ln142_56_fu_6808_p1 = $signed(threshs_m_thresholds_224_q0);

assign sext_ln142_57_fu_7829_p1 = $signed(threshs_m_thresholds_150_q0);

assign sext_ln142_58_fu_7848_p1 = $signed(threshs_m_thresholds_149_q0);

assign sext_ln142_59_fu_7867_p1 = $signed(threshs_m_thresholds_148_q0);

assign sext_ln142_5_fu_4677_p1 = $signed(threshs_m_thresholds_97_q0);

assign sext_ln142_60_fu_7886_p1 = $signed(threshs_m_thresholds_147_q0);

assign sext_ln142_61_fu_7905_p1 = $signed(threshs_m_thresholds_146_q0);

assign sext_ln142_62_fu_7924_p1 = $signed(threshs_m_thresholds_145_q0);

assign sext_ln142_63_fu_7943_p1 = $signed(threshs_m_thresholds_144_q0);

assign sext_ln142_64_fu_7962_p1 = $signed(threshs_m_thresholds_143_q0);

assign sext_ln142_65_fu_7981_p1 = $signed(threshs_m_thresholds_140_q0);

assign sext_ln142_66_fu_8000_p1 = $signed(threshs_m_thresholds_139_q0);

assign sext_ln142_67_fu_8019_p1 = $signed(threshs_m_thresholds_138_q0);

assign sext_ln142_68_fu_8038_p1 = $signed(threshs_m_thresholds_137_q0);

assign sext_ln142_69_fu_8057_p1 = $signed(threshs_m_thresholds_136_q0);

assign sext_ln142_6_fu_4700_p1 = $signed(threshs_m_thresholds_86_q0);

assign sext_ln142_70_fu_8076_p1 = $signed(threshs_m_thresholds_135_q0);

assign sext_ln142_71_fu_8095_p1 = $signed(threshs_m_thresholds_134_q0);

assign sext_ln142_72_fu_8114_p1 = $signed(threshs_m_thresholds_133_q0);

assign sext_ln142_73_fu_8133_p1 = $signed(threshs_m_thresholds_132_q0);

assign sext_ln142_74_fu_8152_p1 = $signed(threshs_m_thresholds_131_q0);

assign sext_ln142_75_fu_8171_p1 = $signed(threshs_m_thresholds_129_q0);

assign sext_ln142_76_fu_8190_p1 = $signed(threshs_m_thresholds_128_q0);

assign sext_ln142_77_fu_8209_p1 = $signed(threshs_m_thresholds_127_q0);

assign sext_ln142_78_fu_8228_p1 = $signed(threshs_m_thresholds_126_q0);

assign sext_ln142_79_fu_8247_p1 = $signed(threshs_m_thresholds_125_q0);

assign sext_ln142_7_fu_4723_p1 = $signed(threshs_m_thresholds_80_q0);

assign sext_ln142_80_fu_8266_p1 = $signed(threshs_m_thresholds_124_q0);

assign sext_ln142_81_fu_8285_p1 = $signed(threshs_m_thresholds_123_q0);

assign sext_ln142_82_fu_8304_p1 = $signed(threshs_m_thresholds_122_q0);

assign sext_ln142_83_fu_8323_p1 = $signed(threshs_m_thresholds_121_q0);

assign sext_ln142_84_fu_8342_p1 = $signed(threshs_m_thresholds_120_q0);

assign sext_ln142_85_fu_8361_p1 = $signed(threshs_m_thresholds_118_q0);

assign sext_ln142_86_fu_8380_p1 = $signed(threshs_m_thresholds_117_q0);

assign sext_ln142_87_fu_8399_p1 = $signed(threshs_m_thresholds_116_q0);

assign sext_ln142_88_fu_8418_p1 = $signed(threshs_m_thresholds_115_q0);

assign sext_ln142_89_fu_8437_p1 = $signed(threshs_m_thresholds_114_q0);

assign sext_ln142_8_fu_4746_p1 = $signed(threshs_m_thresholds_79_q0);

assign sext_ln142_90_fu_8456_p1 = $signed(threshs_m_thresholds_113_q0);

assign sext_ln142_91_fu_8475_p1 = $signed(threshs_m_thresholds_112_q0);

assign sext_ln142_92_fu_8494_p1 = $signed(threshs_m_thresholds_111_q0);

assign sext_ln142_93_fu_8513_p1 = $signed(threshs_m_thresholds_110_q0);

assign sext_ln142_94_fu_8532_p1 = $signed(threshs_m_thresholds_109_q0);

assign sext_ln142_95_fu_8551_p1 = $signed(threshs_m_thresholds_107_q0);

assign sext_ln142_96_fu_8570_p1 = $signed(threshs_m_thresholds_106_q0);

assign sext_ln142_97_fu_8589_p1 = $signed(threshs_m_thresholds_105_q0);

assign sext_ln142_98_fu_8608_p1 = $signed(threshs_m_thresholds_104_q0);

assign sext_ln142_99_fu_8627_p1 = $signed(threshs_m_thresholds_103_q0);

assign sext_ln142_9_fu_4769_p1 = $signed(threshs_m_thresholds_78_q0);

assign sext_ln142_fu_4288_p1 = $signed(threshs_m_thresholds_54_q0);

assign threshs_m_thresholds_100_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_101_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_102_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_103_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_104_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_105_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_106_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_107_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_108_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_109_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_10_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_110_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_111_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_112_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_113_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_114_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_115_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_116_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_117_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_118_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_119_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_11_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_120_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_121_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_122_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_123_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_124_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_125_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_126_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_127_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_128_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_129_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_12_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_130_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_131_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_132_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_133_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_134_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_135_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_136_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_137_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_138_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_139_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_13_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_140_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_141_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_142_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_143_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_144_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_145_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_146_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_147_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_148_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_149_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_14_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_150_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_151_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_152_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_153_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_154_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_155_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_156_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_157_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_158_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_159_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_15_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_160_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_161_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_162_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_163_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_164_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_165_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_166_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_167_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_168_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_169_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_16_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_170_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_171_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_172_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_173_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_174_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_175_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_176_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_177_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_178_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_179_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_17_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_180_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_181_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_182_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_183_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_184_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_185_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_186_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_187_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_188_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_189_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_18_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_190_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_191_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_192_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_193_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_194_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_195_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_196_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_197_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_198_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_199_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_19_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_1_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_200_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_201_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_202_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_203_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_204_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_205_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_206_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_207_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_208_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_209_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_20_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_210_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_211_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_212_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_213_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_214_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_215_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_216_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_217_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_218_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_219_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_21_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_220_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_221_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_222_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_223_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_224_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_225_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_226_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_227_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_228_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_229_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_22_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_230_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_231_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_232_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_233_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_234_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_235_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_236_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_237_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_238_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_239_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_23_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_240_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_241_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_242_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_243_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_244_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_245_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_246_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_247_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_248_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_249_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_24_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_250_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_251_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_252_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_253_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_254_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_25_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_26_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_27_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_28_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_29_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_2_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_30_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_31_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_32_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_33_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_34_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_35_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_36_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_37_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_38_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_39_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_3_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_40_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_41_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_42_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_43_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_44_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_45_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_46_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_47_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_48_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_49_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_4_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_50_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_51_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_52_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_53_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_54_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_55_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_56_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_57_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_58_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_59_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_5_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_60_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_61_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_62_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_63_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_64_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_65_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_66_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_67_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_68_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_69_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_6_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_70_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_71_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_72_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_73_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_74_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_75_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_76_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_77_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_78_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_79_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_7_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_80_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_81_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_82_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_83_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_84_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_85_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_86_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_87_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_88_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_89_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_8_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_90_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_91_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_92_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_93_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_94_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_95_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_96_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_97_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_98_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_99_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_9_address0 = zext_ln142_fu_3940_p1;

assign threshs_m_thresholds_address0 = zext_ln142_fu_3940_p1;

assign xor_ln899_100_fu_6246_p2 = (icmp_ln899_100_fu_6241_p2 ^ 1'd1);

assign xor_ln899_101_fu_6269_p2 = (icmp_ln899_101_fu_6264_p2 ^ 1'd1);

assign xor_ln899_102_fu_6292_p2 = (icmp_ln899_102_fu_6287_p2 ^ 1'd1);

assign xor_ln899_103_fu_6315_p2 = (icmp_ln899_103_fu_6310_p2 ^ 1'd1);

assign xor_ln899_104_fu_6338_p2 = (icmp_ln899_104_fu_6333_p2 ^ 1'd1);

assign xor_ln899_105_fu_6361_p2 = (icmp_ln899_105_fu_6356_p2 ^ 1'd1);

assign xor_ln899_106_fu_6384_p2 = (icmp_ln899_106_fu_6379_p2 ^ 1'd1);

assign xor_ln899_107_fu_6407_p2 = (icmp_ln899_107_fu_6402_p2 ^ 1'd1);

assign xor_ln899_108_fu_6430_p2 = (icmp_ln899_108_fu_6425_p2 ^ 1'd1);

assign xor_ln899_109_fu_6453_p2 = (icmp_ln899_109_fu_6448_p2 ^ 1'd1);

assign xor_ln899_10_fu_4400_p2 = (icmp_ln899_10_fu_4395_p2 ^ 1'd1);

assign xor_ln899_110_fu_6476_p2 = (icmp_ln899_110_fu_6471_p2 ^ 1'd1);

assign xor_ln899_111_fu_6499_p2 = (icmp_ln899_111_fu_6494_p2 ^ 1'd1);

assign xor_ln899_112_fu_6522_p2 = (icmp_ln899_112_fu_6517_p2 ^ 1'd1);

assign xor_ln899_113_fu_6545_p2 = (icmp_ln899_113_fu_6540_p2 ^ 1'd1);

assign xor_ln899_114_fu_6568_p2 = (icmp_ln899_114_fu_6563_p2 ^ 1'd1);

assign xor_ln899_115_fu_6591_p2 = (icmp_ln899_115_fu_6586_p2 ^ 1'd1);

assign xor_ln899_116_fu_6614_p2 = (icmp_ln899_116_fu_6609_p2 ^ 1'd1);

assign xor_ln899_117_fu_6637_p2 = (icmp_ln899_117_fu_6632_p2 ^ 1'd1);

assign xor_ln899_118_fu_6660_p2 = (icmp_ln899_118_fu_6655_p2 ^ 1'd1);

assign xor_ln899_119_fu_6683_p2 = (icmp_ln899_119_fu_6678_p2 ^ 1'd1);

assign xor_ln899_11_fu_4423_p2 = (icmp_ln899_11_fu_4418_p2 ^ 1'd1);

assign xor_ln899_120_fu_6706_p2 = (icmp_ln899_120_fu_6701_p2 ^ 1'd1);

assign xor_ln899_121_fu_6729_p2 = (icmp_ln899_121_fu_6724_p2 ^ 1'd1);

assign xor_ln899_122_fu_6752_p2 = (icmp_ln899_122_fu_6747_p2 ^ 1'd1);

assign xor_ln899_123_fu_6775_p2 = (icmp_ln899_123_fu_6770_p2 ^ 1'd1);

assign xor_ln899_124_fu_6798_p2 = (icmp_ln899_124_fu_6793_p2 ^ 1'd1);

assign xor_ln899_125_fu_6821_p2 = (icmp_ln899_125_fu_6816_p2 ^ 1'd1);

assign xor_ln899_126_fu_6844_p2 = (icmp_ln899_126_fu_6839_p2 ^ 1'd1);

assign xor_ln899_127_fu_6859_p2 = (icmp_ln899_127_fu_6854_p2 ^ 1'd1);

assign xor_ln899_128_fu_6874_p2 = (icmp_ln899_128_fu_6869_p2 ^ 1'd1);

assign xor_ln899_129_fu_6889_p2 = (icmp_ln899_129_fu_6884_p2 ^ 1'd1);

assign xor_ln899_12_fu_4446_p2 = (icmp_ln899_12_fu_4441_p2 ^ 1'd1);

assign xor_ln899_130_fu_6904_p2 = (icmp_ln899_130_fu_6899_p2 ^ 1'd1);

assign xor_ln899_131_fu_6919_p2 = (icmp_ln899_131_fu_6914_p2 ^ 1'd1);

assign xor_ln899_132_fu_6934_p2 = (icmp_ln899_132_fu_6929_p2 ^ 1'd1);

assign xor_ln899_133_fu_6949_p2 = (icmp_ln899_133_fu_6944_p2 ^ 1'd1);

assign xor_ln899_134_fu_6964_p2 = (icmp_ln899_134_fu_6959_p2 ^ 1'd1);

assign xor_ln899_135_fu_6979_p2 = (icmp_ln899_135_fu_6974_p2 ^ 1'd1);

assign xor_ln899_136_fu_6994_p2 = (icmp_ln899_136_fu_6989_p2 ^ 1'd1);

assign xor_ln899_137_fu_7009_p2 = (icmp_ln899_137_fu_7004_p2 ^ 1'd1);

assign xor_ln899_138_fu_7024_p2 = (icmp_ln899_138_fu_7019_p2 ^ 1'd1);

assign xor_ln899_139_fu_7039_p2 = (icmp_ln899_139_fu_7034_p2 ^ 1'd1);

assign xor_ln899_13_fu_4469_p2 = (icmp_ln899_13_fu_4464_p2 ^ 1'd1);

assign xor_ln899_140_fu_7054_p2 = (icmp_ln899_140_fu_7049_p2 ^ 1'd1);

assign xor_ln899_141_fu_7069_p2 = (icmp_ln899_141_fu_7064_p2 ^ 1'd1);

assign xor_ln899_142_fu_7084_p2 = (icmp_ln899_142_fu_7079_p2 ^ 1'd1);

assign xor_ln899_143_fu_7099_p2 = (icmp_ln899_143_fu_7094_p2 ^ 1'd1);

assign xor_ln899_144_fu_7114_p2 = (icmp_ln899_144_fu_7109_p2 ^ 1'd1);

assign xor_ln899_145_fu_7129_p2 = (icmp_ln899_145_fu_7124_p2 ^ 1'd1);

assign xor_ln899_146_fu_7144_p2 = (icmp_ln899_146_fu_7139_p2 ^ 1'd1);

assign xor_ln899_147_fu_7159_p2 = (icmp_ln899_147_fu_7154_p2 ^ 1'd1);

assign xor_ln899_148_fu_7174_p2 = (icmp_ln899_148_fu_7169_p2 ^ 1'd1);

assign xor_ln899_149_fu_7189_p2 = (icmp_ln899_149_fu_7184_p2 ^ 1'd1);

assign xor_ln899_14_fu_4492_p2 = (icmp_ln899_14_fu_4487_p2 ^ 1'd1);

assign xor_ln899_150_fu_7204_p2 = (icmp_ln899_150_fu_7199_p2 ^ 1'd1);

assign xor_ln899_151_fu_7219_p2 = (icmp_ln899_151_fu_7214_p2 ^ 1'd1);

assign xor_ln899_152_fu_7234_p2 = (icmp_ln899_152_fu_7229_p2 ^ 1'd1);

assign xor_ln899_153_fu_7249_p2 = (icmp_ln899_153_fu_7244_p2 ^ 1'd1);

assign xor_ln899_154_fu_7264_p2 = (icmp_ln899_154_fu_7259_p2 ^ 1'd1);

assign xor_ln899_155_fu_7279_p2 = (icmp_ln899_155_fu_7274_p2 ^ 1'd1);

assign xor_ln899_156_fu_7294_p2 = (icmp_ln899_156_fu_7289_p2 ^ 1'd1);

assign xor_ln899_157_fu_7309_p2 = (icmp_ln899_157_fu_7304_p2 ^ 1'd1);

assign xor_ln899_158_fu_7324_p2 = (icmp_ln899_158_fu_7319_p2 ^ 1'd1);

assign xor_ln899_159_fu_7339_p2 = (icmp_ln899_159_fu_7334_p2 ^ 1'd1);

assign xor_ln899_15_fu_4511_p2 = (icmp_ln899_15_fu_4506_p2 ^ 1'd1);

assign xor_ln899_160_fu_7354_p2 = (icmp_ln899_160_fu_7349_p2 ^ 1'd1);

assign xor_ln899_161_fu_7369_p2 = (icmp_ln899_161_fu_7364_p2 ^ 1'd1);

assign xor_ln899_162_fu_7384_p2 = (icmp_ln899_162_fu_7379_p2 ^ 1'd1);

assign xor_ln899_163_fu_7399_p2 = (icmp_ln899_163_fu_7394_p2 ^ 1'd1);

assign xor_ln899_164_fu_7414_p2 = (icmp_ln899_164_fu_7409_p2 ^ 1'd1);

assign xor_ln899_165_fu_7429_p2 = (icmp_ln899_165_fu_7424_p2 ^ 1'd1);

assign xor_ln899_166_fu_7444_p2 = (icmp_ln899_166_fu_7439_p2 ^ 1'd1);

assign xor_ln899_167_fu_7459_p2 = (icmp_ln899_167_fu_7454_p2 ^ 1'd1);

assign xor_ln899_168_fu_7474_p2 = (icmp_ln899_168_fu_7469_p2 ^ 1'd1);

assign xor_ln899_169_fu_7489_p2 = (icmp_ln899_169_fu_7484_p2 ^ 1'd1);

assign xor_ln899_16_fu_4530_p2 = (icmp_ln899_16_fu_4525_p2 ^ 1'd1);

assign xor_ln899_170_fu_7504_p2 = (icmp_ln899_170_fu_7499_p2 ^ 1'd1);

assign xor_ln899_171_fu_7519_p2 = (icmp_ln899_171_fu_7514_p2 ^ 1'd1);

assign xor_ln899_172_fu_7534_p2 = (icmp_ln899_172_fu_7529_p2 ^ 1'd1);

assign xor_ln899_173_fu_7549_p2 = (icmp_ln899_173_fu_7544_p2 ^ 1'd1);

assign xor_ln899_174_fu_7564_p2 = (icmp_ln899_174_fu_7559_p2 ^ 1'd1);

assign xor_ln899_175_fu_7579_p2 = (icmp_ln899_175_fu_7574_p2 ^ 1'd1);

assign xor_ln899_176_fu_7594_p2 = (icmp_ln899_176_fu_7589_p2 ^ 1'd1);

assign xor_ln899_177_fu_7609_p2 = (icmp_ln899_177_fu_7604_p2 ^ 1'd1);

assign xor_ln899_178_fu_7624_p2 = (icmp_ln899_178_fu_7619_p2 ^ 1'd1);

assign xor_ln899_179_fu_7639_p2 = (icmp_ln899_179_fu_7634_p2 ^ 1'd1);

assign xor_ln899_17_fu_4549_p2 = (icmp_ln899_17_fu_4544_p2 ^ 1'd1);

assign xor_ln899_180_fu_7654_p2 = (icmp_ln899_180_fu_7649_p2 ^ 1'd1);

assign xor_ln899_181_fu_7669_p2 = (icmp_ln899_181_fu_7664_p2 ^ 1'd1);

assign xor_ln899_182_fu_7684_p2 = (icmp_ln899_182_fu_7679_p2 ^ 1'd1);

assign xor_ln899_183_fu_7699_p2 = (icmp_ln899_183_fu_7694_p2 ^ 1'd1);

assign xor_ln899_184_fu_7714_p2 = (icmp_ln899_184_fu_7709_p2 ^ 1'd1);

assign xor_ln899_185_fu_7729_p2 = (icmp_ln899_185_fu_7724_p2 ^ 1'd1);

assign xor_ln899_186_fu_7744_p2 = (icmp_ln899_186_fu_7739_p2 ^ 1'd1);

assign xor_ln899_187_fu_7759_p2 = (icmp_ln899_187_fu_7754_p2 ^ 1'd1);

assign xor_ln899_188_fu_7774_p2 = (icmp_ln899_188_fu_7769_p2 ^ 1'd1);

assign xor_ln899_189_fu_7789_p2 = (icmp_ln899_189_fu_7784_p2 ^ 1'd1);

assign xor_ln899_18_fu_4568_p2 = (icmp_ln899_18_fu_4563_p2 ^ 1'd1);

assign xor_ln899_190_fu_7804_p2 = (icmp_ln899_190_fu_7799_p2 ^ 1'd1);

assign xor_ln899_191_fu_7819_p2 = (icmp_ln899_191_fu_7814_p2 ^ 1'd1);

assign xor_ln899_192_fu_7838_p2 = (icmp_ln899_192_fu_7833_p2 ^ 1'd1);

assign xor_ln899_193_fu_7857_p2 = (icmp_ln899_193_fu_7852_p2 ^ 1'd1);

assign xor_ln899_194_fu_7876_p2 = (icmp_ln899_194_fu_7871_p2 ^ 1'd1);

assign xor_ln899_195_fu_7895_p2 = (icmp_ln899_195_fu_7890_p2 ^ 1'd1);

assign xor_ln899_196_fu_7914_p2 = (icmp_ln899_196_fu_7909_p2 ^ 1'd1);

assign xor_ln899_197_fu_7933_p2 = (icmp_ln899_197_fu_7928_p2 ^ 1'd1);

assign xor_ln899_198_fu_7952_p2 = (icmp_ln899_198_fu_7947_p2 ^ 1'd1);

assign xor_ln899_199_fu_7971_p2 = (icmp_ln899_199_fu_7966_p2 ^ 1'd1);

assign xor_ln899_19_fu_4587_p2 = (icmp_ln899_19_fu_4582_p2 ^ 1'd1);

assign xor_ln899_1_fu_10677_p2 = (icmp_ln899_1_reg_13050 ^ 1'd1);

assign xor_ln899_200_fu_7990_p2 = (icmp_ln899_200_fu_7985_p2 ^ 1'd1);

assign xor_ln899_201_fu_8009_p2 = (icmp_ln899_201_fu_8004_p2 ^ 1'd1);

assign xor_ln899_202_fu_8028_p2 = (icmp_ln899_202_fu_8023_p2 ^ 1'd1);

assign xor_ln899_203_fu_8047_p2 = (icmp_ln899_203_fu_8042_p2 ^ 1'd1);

assign xor_ln899_204_fu_8066_p2 = (icmp_ln899_204_fu_8061_p2 ^ 1'd1);

assign xor_ln899_205_fu_8085_p2 = (icmp_ln899_205_fu_8080_p2 ^ 1'd1);

assign xor_ln899_206_fu_8104_p2 = (icmp_ln899_206_fu_8099_p2 ^ 1'd1);

assign xor_ln899_207_fu_8123_p2 = (icmp_ln899_207_fu_8118_p2 ^ 1'd1);

assign xor_ln899_208_fu_8142_p2 = (icmp_ln899_208_fu_8137_p2 ^ 1'd1);

assign xor_ln899_209_fu_8161_p2 = (icmp_ln899_209_fu_8156_p2 ^ 1'd1);

assign xor_ln899_20_fu_4606_p2 = (icmp_ln899_20_fu_4601_p2 ^ 1'd1);

assign xor_ln899_210_fu_8180_p2 = (icmp_ln899_210_fu_8175_p2 ^ 1'd1);

assign xor_ln899_211_fu_8199_p2 = (icmp_ln899_211_fu_8194_p2 ^ 1'd1);

assign xor_ln899_212_fu_8218_p2 = (icmp_ln899_212_fu_8213_p2 ^ 1'd1);

assign xor_ln899_213_fu_8237_p2 = (icmp_ln899_213_fu_8232_p2 ^ 1'd1);

assign xor_ln899_214_fu_8256_p2 = (icmp_ln899_214_fu_8251_p2 ^ 1'd1);

assign xor_ln899_215_fu_8275_p2 = (icmp_ln899_215_fu_8270_p2 ^ 1'd1);

assign xor_ln899_216_fu_8294_p2 = (icmp_ln899_216_fu_8289_p2 ^ 1'd1);

assign xor_ln899_217_fu_8313_p2 = (icmp_ln899_217_fu_8308_p2 ^ 1'd1);

assign xor_ln899_218_fu_8332_p2 = (icmp_ln899_218_fu_8327_p2 ^ 1'd1);

assign xor_ln899_219_fu_8351_p2 = (icmp_ln899_219_fu_8346_p2 ^ 1'd1);

assign xor_ln899_21_fu_4625_p2 = (icmp_ln899_21_fu_4620_p2 ^ 1'd1);

assign xor_ln899_220_fu_8370_p2 = (icmp_ln899_220_fu_8365_p2 ^ 1'd1);

assign xor_ln899_221_fu_8389_p2 = (icmp_ln899_221_fu_8384_p2 ^ 1'd1);

assign xor_ln899_222_fu_8408_p2 = (icmp_ln899_222_fu_8403_p2 ^ 1'd1);

assign xor_ln899_223_fu_8427_p2 = (icmp_ln899_223_fu_8422_p2 ^ 1'd1);

assign xor_ln899_224_fu_8446_p2 = (icmp_ln899_224_fu_8441_p2 ^ 1'd1);

assign xor_ln899_225_fu_8465_p2 = (icmp_ln899_225_fu_8460_p2 ^ 1'd1);

assign xor_ln899_226_fu_8484_p2 = (icmp_ln899_226_fu_8479_p2 ^ 1'd1);

assign xor_ln899_227_fu_8503_p2 = (icmp_ln899_227_fu_8498_p2 ^ 1'd1);

assign xor_ln899_228_fu_8522_p2 = (icmp_ln899_228_fu_8517_p2 ^ 1'd1);

assign xor_ln899_229_fu_8541_p2 = (icmp_ln899_229_fu_8536_p2 ^ 1'd1);

assign xor_ln899_22_fu_4644_p2 = (icmp_ln899_22_fu_4639_p2 ^ 1'd1);

assign xor_ln899_230_fu_8560_p2 = (icmp_ln899_230_fu_8555_p2 ^ 1'd1);

assign xor_ln899_231_fu_8579_p2 = (icmp_ln899_231_fu_8574_p2 ^ 1'd1);

assign xor_ln899_232_fu_8598_p2 = (icmp_ln899_232_fu_8593_p2 ^ 1'd1);

assign xor_ln899_233_fu_8617_p2 = (icmp_ln899_233_fu_8612_p2 ^ 1'd1);

assign xor_ln899_234_fu_8636_p2 = (icmp_ln899_234_fu_8631_p2 ^ 1'd1);

assign xor_ln899_235_fu_8655_p2 = (icmp_ln899_235_fu_8650_p2 ^ 1'd1);

assign xor_ln899_236_fu_8674_p2 = (icmp_ln899_236_fu_8669_p2 ^ 1'd1);

assign xor_ln899_237_fu_8693_p2 = (icmp_ln899_237_fu_8688_p2 ^ 1'd1);

assign xor_ln899_238_fu_8712_p2 = (icmp_ln899_238_fu_8707_p2 ^ 1'd1);

assign xor_ln899_239_fu_8731_p2 = (icmp_ln899_239_fu_8726_p2 ^ 1'd1);

assign xor_ln899_23_fu_4667_p2 = (icmp_ln899_23_fu_4662_p2 ^ 1'd1);

assign xor_ln899_240_fu_8750_p2 = (icmp_ln899_240_fu_8745_p2 ^ 1'd1);

assign xor_ln899_241_fu_8769_p2 = (icmp_ln899_241_fu_8764_p2 ^ 1'd1);

assign xor_ln899_242_fu_8788_p2 = (icmp_ln899_242_fu_8783_p2 ^ 1'd1);

assign xor_ln899_243_fu_8807_p2 = (icmp_ln899_243_fu_8802_p2 ^ 1'd1);

assign xor_ln899_244_fu_8826_p2 = (icmp_ln899_244_fu_8821_p2 ^ 1'd1);

assign xor_ln899_245_fu_8845_p2 = (icmp_ln899_245_fu_8840_p2 ^ 1'd1);

assign xor_ln899_246_fu_8864_p2 = (icmp_ln899_246_fu_8859_p2 ^ 1'd1);

assign xor_ln899_247_fu_8883_p2 = (icmp_ln899_247_fu_8878_p2 ^ 1'd1);

assign xor_ln899_248_fu_8902_p2 = (icmp_ln899_248_fu_8897_p2 ^ 1'd1);

assign xor_ln899_249_fu_8921_p2 = (icmp_ln899_249_fu_8916_p2 ^ 1'd1);

assign xor_ln899_24_fu_4690_p2 = (icmp_ln899_24_fu_4685_p2 ^ 1'd1);

assign xor_ln899_250_fu_8940_p2 = (icmp_ln899_250_fu_8935_p2 ^ 1'd1);

assign xor_ln899_251_fu_8959_p2 = (icmp_ln899_251_fu_8954_p2 ^ 1'd1);

assign xor_ln899_252_fu_8978_p2 = (icmp_ln899_252_fu_8973_p2 ^ 1'd1);

assign xor_ln899_253_fu_8997_p2 = (icmp_ln899_253_fu_8992_p2 ^ 1'd1);

assign xor_ln899_254_fu_9016_p2 = (icmp_ln899_254_fu_9011_p2 ^ 1'd1);

assign xor_ln899_25_fu_4713_p2 = (icmp_ln899_25_fu_4708_p2 ^ 1'd1);

assign xor_ln899_26_fu_4736_p2 = (icmp_ln899_26_fu_4731_p2 ^ 1'd1);

assign xor_ln899_27_fu_4759_p2 = (icmp_ln899_27_fu_4754_p2 ^ 1'd1);

assign xor_ln899_28_fu_4782_p2 = (icmp_ln899_28_fu_4777_p2 ^ 1'd1);

assign xor_ln899_29_fu_4805_p2 = (icmp_ln899_29_fu_4800_p2 ^ 1'd1);

assign xor_ln899_2_fu_10686_p2 = (icmp_ln899_2_reg_13055 ^ 1'd1);

assign xor_ln899_30_fu_4828_p2 = (icmp_ln899_30_fu_4823_p2 ^ 1'd1);

assign xor_ln899_31_fu_4847_p2 = (icmp_ln899_31_fu_4842_p2 ^ 1'd1);

assign xor_ln899_32_fu_4866_p2 = (icmp_ln899_32_fu_4861_p2 ^ 1'd1);

assign xor_ln899_33_fu_4885_p2 = (icmp_ln899_33_fu_4880_p2 ^ 1'd1);

assign xor_ln899_34_fu_4904_p2 = (icmp_ln899_34_fu_4899_p2 ^ 1'd1);

assign xor_ln899_35_fu_4923_p2 = (icmp_ln899_35_fu_4918_p2 ^ 1'd1);

assign xor_ln899_36_fu_4942_p2 = (icmp_ln899_36_fu_4937_p2 ^ 1'd1);

assign xor_ln899_37_fu_4961_p2 = (icmp_ln899_37_fu_4956_p2 ^ 1'd1);

assign xor_ln899_38_fu_4980_p2 = (icmp_ln899_38_fu_4975_p2 ^ 1'd1);

assign xor_ln899_39_fu_4999_p2 = (icmp_ln899_39_fu_4994_p2 ^ 1'd1);

assign xor_ln899_3_fu_4259_p2 = (icmp_ln899_3_fu_4254_p2 ^ 1'd1);

assign xor_ln899_40_fu_5018_p2 = (icmp_ln899_40_fu_5013_p2 ^ 1'd1);

assign xor_ln899_41_fu_5037_p2 = (icmp_ln899_41_fu_5032_p2 ^ 1'd1);

assign xor_ln899_42_fu_5056_p2 = (icmp_ln899_42_fu_5051_p2 ^ 1'd1);

assign xor_ln899_43_fu_5075_p2 = (icmp_ln899_43_fu_5070_p2 ^ 1'd1);

assign xor_ln899_44_fu_5094_p2 = (icmp_ln899_44_fu_5089_p2 ^ 1'd1);

assign xor_ln899_45_fu_5113_p2 = (icmp_ln899_45_fu_5108_p2 ^ 1'd1);

assign xor_ln899_46_fu_5132_p2 = (icmp_ln899_46_fu_5127_p2 ^ 1'd1);

assign xor_ln899_47_fu_5155_p2 = (icmp_ln899_47_fu_5150_p2 ^ 1'd1);

assign xor_ln899_48_fu_5178_p2 = (icmp_ln899_48_fu_5173_p2 ^ 1'd1);

assign xor_ln899_49_fu_5201_p2 = (icmp_ln899_49_fu_5196_p2 ^ 1'd1);

assign xor_ln899_4_fu_4278_p2 = (icmp_ln899_4_fu_4273_p2 ^ 1'd1);

assign xor_ln899_50_fu_5224_p2 = (icmp_ln899_50_fu_5219_p2 ^ 1'd1);

assign xor_ln899_51_fu_5247_p2 = (icmp_ln899_51_fu_5242_p2 ^ 1'd1);

assign xor_ln899_52_fu_5270_p2 = (icmp_ln899_52_fu_5265_p2 ^ 1'd1);

assign xor_ln899_53_fu_5293_p2 = (icmp_ln899_53_fu_5288_p2 ^ 1'd1);

assign xor_ln899_54_fu_5316_p2 = (icmp_ln899_54_fu_5311_p2 ^ 1'd1);

assign xor_ln899_55_fu_5339_p2 = (icmp_ln899_55_fu_5334_p2 ^ 1'd1);

assign xor_ln899_56_fu_5362_p2 = (icmp_ln899_56_fu_5357_p2 ^ 1'd1);

assign xor_ln899_57_fu_5385_p2 = (icmp_ln899_57_fu_5380_p2 ^ 1'd1);

assign xor_ln899_58_fu_5408_p2 = (icmp_ln899_58_fu_5403_p2 ^ 1'd1);

assign xor_ln899_59_fu_5431_p2 = (icmp_ln899_59_fu_5426_p2 ^ 1'd1);

assign xor_ln899_5_fu_4301_p2 = (icmp_ln899_5_fu_4296_p2 ^ 1'd1);

assign xor_ln899_60_fu_5454_p2 = (icmp_ln899_60_fu_5449_p2 ^ 1'd1);

assign xor_ln899_61_fu_5477_p2 = (icmp_ln899_61_fu_5472_p2 ^ 1'd1);

assign xor_ln899_62_fu_5500_p2 = (icmp_ln899_62_fu_5495_p2 ^ 1'd1);

assign xor_ln899_63_fu_5519_p2 = (icmp_ln899_63_fu_5514_p2 ^ 1'd1);

assign xor_ln899_64_fu_5538_p2 = (icmp_ln899_64_fu_5533_p2 ^ 1'd1);

assign xor_ln899_65_fu_5557_p2 = (icmp_ln899_65_fu_5552_p2 ^ 1'd1);

assign xor_ln899_66_fu_5576_p2 = (icmp_ln899_66_fu_5571_p2 ^ 1'd1);

assign xor_ln899_67_fu_5595_p2 = (icmp_ln899_67_fu_5590_p2 ^ 1'd1);

assign xor_ln899_68_fu_5614_p2 = (icmp_ln899_68_fu_5609_p2 ^ 1'd1);

assign xor_ln899_69_fu_5633_p2 = (icmp_ln899_69_fu_5628_p2 ^ 1'd1);

assign xor_ln899_6_fu_4324_p2 = (icmp_ln899_6_fu_4319_p2 ^ 1'd1);

assign xor_ln899_70_fu_5652_p2 = (icmp_ln899_70_fu_5647_p2 ^ 1'd1);

assign xor_ln899_71_fu_5671_p2 = (icmp_ln899_71_fu_5666_p2 ^ 1'd1);

assign xor_ln899_72_fu_5690_p2 = (icmp_ln899_72_fu_5685_p2 ^ 1'd1);

assign xor_ln899_73_fu_5709_p2 = (icmp_ln899_73_fu_5704_p2 ^ 1'd1);

assign xor_ln899_74_fu_5728_p2 = (icmp_ln899_74_fu_5723_p2 ^ 1'd1);

assign xor_ln899_75_fu_5747_p2 = (icmp_ln899_75_fu_5742_p2 ^ 1'd1);

assign xor_ln899_76_fu_5766_p2 = (icmp_ln899_76_fu_5761_p2 ^ 1'd1);

assign xor_ln899_77_fu_5785_p2 = (icmp_ln899_77_fu_5780_p2 ^ 1'd1);

assign xor_ln899_78_fu_5804_p2 = (icmp_ln899_78_fu_5799_p2 ^ 1'd1);

assign xor_ln899_79_fu_5823_p2 = (icmp_ln899_79_fu_5818_p2 ^ 1'd1);

assign xor_ln899_7_fu_4343_p2 = (icmp_ln899_7_fu_4338_p2 ^ 1'd1);

assign xor_ln899_80_fu_5842_p2 = (icmp_ln899_80_fu_5837_p2 ^ 1'd1);

assign xor_ln899_81_fu_5861_p2 = (icmp_ln899_81_fu_5856_p2 ^ 1'd1);

assign xor_ln899_82_fu_5880_p2 = (icmp_ln899_82_fu_5875_p2 ^ 1'd1);

assign xor_ln899_83_fu_5899_p2 = (icmp_ln899_83_fu_5894_p2 ^ 1'd1);

assign xor_ln899_84_fu_5918_p2 = (icmp_ln899_84_fu_5913_p2 ^ 1'd1);

assign xor_ln899_85_fu_5937_p2 = (icmp_ln899_85_fu_5932_p2 ^ 1'd1);

assign xor_ln899_86_fu_5956_p2 = (icmp_ln899_86_fu_5951_p2 ^ 1'd1);

assign xor_ln899_87_fu_5975_p2 = (icmp_ln899_87_fu_5970_p2 ^ 1'd1);

assign xor_ln899_88_fu_5994_p2 = (icmp_ln899_88_fu_5989_p2 ^ 1'd1);

assign xor_ln899_89_fu_6013_p2 = (icmp_ln899_89_fu_6008_p2 ^ 1'd1);

assign xor_ln899_8_fu_4362_p2 = (icmp_ln899_8_fu_4357_p2 ^ 1'd1);

assign xor_ln899_90_fu_6032_p2 = (icmp_ln899_90_fu_6027_p2 ^ 1'd1);

assign xor_ln899_91_fu_6051_p2 = (icmp_ln899_91_fu_6046_p2 ^ 1'd1);

assign xor_ln899_92_fu_6070_p2 = (icmp_ln899_92_fu_6065_p2 ^ 1'd1);

assign xor_ln899_93_fu_6089_p2 = (icmp_ln899_93_fu_6084_p2 ^ 1'd1);

assign xor_ln899_94_fu_6108_p2 = (icmp_ln899_94_fu_6103_p2 ^ 1'd1);

assign xor_ln899_95_fu_6131_p2 = (icmp_ln899_95_fu_6126_p2 ^ 1'd1);

assign xor_ln899_96_fu_6154_p2 = (icmp_ln899_96_fu_6149_p2 ^ 1'd1);

assign xor_ln899_97_fu_6177_p2 = (icmp_ln899_97_fu_6172_p2 ^ 1'd1);

assign xor_ln899_98_fu_6200_p2 = (icmp_ln899_98_fu_6195_p2 ^ 1'd1);

assign xor_ln899_99_fu_6223_p2 = (icmp_ln899_99_fu_6218_p2 ^ 1'd1);

assign xor_ln899_9_fu_4381_p2 = (icmp_ln899_9_fu_4376_p2 ^ 1'd1);

assign xor_ln899_fu_10664_p2 = (icmp_ln899_reg_13045 ^ 1'd1);

assign zext_ln142_100_fu_5261_p1 = $unsigned(sext_ln142_16_fu_5257_p1);

assign zext_ln142_101_fu_5276_p1 = xor_ln899_52_fu_5270_p2;

assign zext_ln142_102_fu_5284_p1 = $unsigned(sext_ln142_17_fu_5280_p1);

assign zext_ln142_103_fu_5299_p1 = xor_ln899_53_fu_5293_p2;

assign zext_ln142_104_fu_5307_p1 = $unsigned(sext_ln142_18_fu_5303_p1);

assign zext_ln142_105_fu_5322_p1 = xor_ln899_54_fu_5316_p2;

assign zext_ln142_106_fu_5330_p1 = $unsigned(sext_ln142_19_fu_5326_p1);

assign zext_ln142_107_fu_5345_p1 = xor_ln899_55_fu_5339_p2;

assign zext_ln142_108_fu_5353_p1 = $unsigned(sext_ln142_20_fu_5349_p1);

assign zext_ln142_109_fu_5368_p1 = xor_ln899_56_fu_5362_p2;

assign zext_ln142_10_fu_4307_p1 = xor_ln899_5_fu_4301_p2;

assign zext_ln142_110_fu_5376_p1 = $unsigned(sext_ln142_21_fu_5372_p1);

assign zext_ln142_111_fu_5391_p1 = xor_ln899_57_fu_5385_p2;

assign zext_ln142_112_fu_5399_p1 = $unsigned(sext_ln142_22_fu_5395_p1);

assign zext_ln142_113_fu_5414_p1 = xor_ln899_58_fu_5408_p2;

assign zext_ln142_114_fu_5422_p1 = $unsigned(sext_ln142_23_fu_5418_p1);

assign zext_ln142_115_fu_5437_p1 = xor_ln899_59_fu_5431_p2;

assign zext_ln142_116_fu_5445_p1 = $unsigned(sext_ln142_24_fu_5441_p1);

assign zext_ln142_117_fu_5460_p1 = xor_ln899_60_fu_5454_p2;

assign zext_ln142_118_fu_5468_p1 = $unsigned(sext_ln142_25_fu_5464_p1);

assign zext_ln142_119_fu_5483_p1 = xor_ln899_61_fu_5477_p2;

assign zext_ln142_11_fu_4330_p1 = xor_ln899_6_fu_4324_p2;

assign zext_ln142_120_fu_5506_p1 = xor_ln899_62_fu_5500_p2;

assign zext_ln142_121_fu_5510_p1 = threshs_m_thresholds_39_q0;

assign zext_ln142_122_fu_5525_p1 = xor_ln899_63_fu_5519_p2;

assign zext_ln142_123_fu_5529_p1 = threshs_m_thresholds_38_q0;

assign zext_ln142_124_fu_5544_p1 = xor_ln899_64_fu_5538_p2;

assign zext_ln142_125_fu_5548_p1 = threshs_m_thresholds_37_q0;

assign zext_ln142_126_fu_5563_p1 = xor_ln899_65_fu_5557_p2;

assign zext_ln142_127_fu_5567_p1 = threshs_m_thresholds_36_q0;

assign zext_ln142_128_fu_5582_p1 = xor_ln899_66_fu_5576_p2;

assign zext_ln142_129_fu_5586_p1 = threshs_m_thresholds_35_q0;

assign zext_ln142_12_fu_4334_p1 = threshs_m_thresholds_32_q0;

assign zext_ln142_130_fu_5601_p1 = xor_ln899_67_fu_5595_p2;

assign zext_ln142_131_fu_5605_p1 = threshs_m_thresholds_34_q0;

assign zext_ln142_132_fu_5620_p1 = xor_ln899_68_fu_5614_p2;

assign zext_ln142_133_fu_5624_p1 = threshs_m_thresholds_33_q0;

assign zext_ln142_134_fu_5639_p1 = xor_ln899_69_fu_5633_p2;

assign zext_ln142_135_fu_5643_p1 = threshs_m_thresholds_31_q0;

assign zext_ln142_136_fu_5658_p1 = xor_ln899_70_fu_5652_p2;

assign zext_ln142_137_fu_5662_p1 = threshs_m_thresholds_30_q0;

assign zext_ln142_138_fu_5677_p1 = xor_ln899_71_fu_5671_p2;

assign zext_ln142_139_fu_5681_p1 = threshs_m_thresholds_29_q0;

assign zext_ln142_13_fu_4349_p1 = xor_ln899_7_fu_4343_p2;

assign zext_ln142_140_fu_5696_p1 = xor_ln899_72_fu_5690_p2;

assign zext_ln142_141_fu_5700_p1 = threshs_m_thresholds_28_q0;

assign zext_ln142_142_fu_5715_p1 = xor_ln899_73_fu_5709_p2;

assign zext_ln142_143_fu_5719_p1 = threshs_m_thresholds_27_q0;

assign zext_ln142_144_fu_5734_p1 = xor_ln899_74_fu_5728_p2;

assign zext_ln142_145_fu_5738_p1 = threshs_m_thresholds_26_q0;

assign zext_ln142_146_fu_5753_p1 = xor_ln899_75_fu_5747_p2;

assign zext_ln142_147_fu_5757_p1 = threshs_m_thresholds_25_q0;

assign zext_ln142_148_fu_5772_p1 = xor_ln899_76_fu_5766_p2;

assign zext_ln142_149_fu_5776_p1 = threshs_m_thresholds_24_q0;

assign zext_ln142_14_fu_4353_p1 = threshs_m_thresholds_21_q0;

assign zext_ln142_150_fu_5791_p1 = xor_ln899_77_fu_5785_p2;

assign zext_ln142_151_fu_5795_p1 = threshs_m_thresholds_23_q0;

assign zext_ln142_152_fu_5810_p1 = xor_ln899_78_fu_5804_p2;

assign zext_ln142_153_fu_5814_p1 = threshs_m_thresholds_22_q0;

assign zext_ln142_154_fu_5829_p1 = xor_ln899_79_fu_5823_p2;

assign zext_ln142_155_fu_5833_p1 = threshs_m_thresholds_20_q0;

assign zext_ln142_156_fu_5848_p1 = xor_ln899_80_fu_5842_p2;

assign zext_ln142_157_fu_5852_p1 = threshs_m_thresholds_19_q0;

assign zext_ln142_158_fu_5867_p1 = xor_ln899_81_fu_5861_p2;

assign zext_ln142_159_fu_5871_p1 = threshs_m_thresholds_18_q0;

assign zext_ln142_15_fu_4368_p1 = xor_ln899_8_fu_4362_p2;

assign zext_ln142_160_fu_5886_p1 = xor_ln899_82_fu_5880_p2;

assign zext_ln142_161_fu_5890_p1 = threshs_m_thresholds_17_q0;

assign zext_ln142_162_fu_5905_p1 = xor_ln899_83_fu_5899_p2;

assign zext_ln142_163_fu_5909_p1 = threshs_m_thresholds_16_q0;

assign zext_ln142_164_fu_5924_p1 = xor_ln899_84_fu_5918_p2;

assign zext_ln142_165_fu_5928_p1 = threshs_m_thresholds_15_q0;

assign zext_ln142_166_fu_5943_p1 = xor_ln899_85_fu_5937_p2;

assign zext_ln142_167_fu_5947_p1 = threshs_m_thresholds_14_q0;

assign zext_ln142_168_fu_5962_p1 = xor_ln899_86_fu_5956_p2;

assign zext_ln142_169_fu_5966_p1 = threshs_m_thresholds_13_q0;

assign zext_ln142_16_fu_4372_p1 = threshs_m_thresholds_10_q0;

assign zext_ln142_170_fu_5981_p1 = xor_ln899_87_fu_5975_p2;

assign zext_ln142_171_fu_5985_p1 = threshs_m_thresholds_12_q0;

assign zext_ln142_172_fu_6000_p1 = xor_ln899_88_fu_5994_p2;

assign zext_ln142_173_fu_6004_p1 = threshs_m_thresholds_11_q0;

assign zext_ln142_174_fu_6019_p1 = xor_ln899_89_fu_6013_p2;

assign zext_ln142_175_fu_6023_p1 = threshs_m_thresholds_9_q0;

assign zext_ln142_176_fu_6038_p1 = xor_ln899_90_fu_6032_p2;

assign zext_ln142_177_fu_6042_p1 = threshs_m_thresholds_8_q0;

assign zext_ln142_178_fu_6057_p1 = xor_ln899_91_fu_6051_p2;

assign zext_ln142_179_fu_6061_p1 = threshs_m_thresholds_7_q0;

assign zext_ln142_17_fu_4387_p1 = xor_ln899_9_fu_4381_p2;

assign zext_ln142_180_fu_6076_p1 = xor_ln899_92_fu_6070_p2;

assign zext_ln142_181_fu_6080_p1 = threshs_m_thresholds_6_q0;

assign zext_ln142_182_fu_6095_p1 = xor_ln899_93_fu_6089_p2;

assign zext_ln142_183_fu_6099_p1 = threshs_m_thresholds_5_q0;

assign zext_ln142_184_fu_6114_p1 = xor_ln899_94_fu_6108_p2;

assign zext_ln142_185_fu_6122_p1 = $unsigned(sext_ln142_26_fu_6118_p1);

assign zext_ln142_186_fu_6137_p1 = xor_ln899_95_fu_6131_p2;

assign zext_ln142_187_fu_6145_p1 = $unsigned(sext_ln142_27_fu_6141_p1);

assign zext_ln142_188_fu_6160_p1 = xor_ln899_96_fu_6154_p2;

assign zext_ln142_189_fu_6168_p1 = $unsigned(sext_ln142_28_fu_6164_p1);

assign zext_ln142_18_fu_4391_p1 = threshs_m_thresholds_252_q0;

assign zext_ln142_190_fu_6183_p1 = xor_ln899_97_fu_6177_p2;

assign zext_ln142_191_fu_6191_p1 = $unsigned(sext_ln142_29_fu_6187_p1);

assign zext_ln142_192_fu_6206_p1 = xor_ln899_98_fu_6200_p2;

assign zext_ln142_193_fu_6214_p1 = $unsigned(sext_ln142_30_fu_6210_p1);

assign zext_ln142_194_fu_6229_p1 = xor_ln899_99_fu_6223_p2;

assign zext_ln142_195_fu_6237_p1 = $unsigned(sext_ln142_31_fu_6233_p1);

assign zext_ln142_196_fu_6252_p1 = xor_ln899_100_fu_6246_p2;

assign zext_ln142_197_fu_6260_p1 = $unsigned(sext_ln142_32_fu_6256_p1);

assign zext_ln142_198_fu_6275_p1 = xor_ln899_101_fu_6269_p2;

assign zext_ln142_199_fu_6283_p1 = $unsigned(sext_ln142_33_fu_6279_p1);

assign zext_ln142_19_fu_4406_p1 = xor_ln899_10_fu_4400_p2;

assign zext_ln142_1_fu_4219_p1 = threshs_m_thresholds_254_q0;

assign zext_ln142_200_fu_6298_p1 = xor_ln899_102_fu_6292_p2;

assign zext_ln142_201_fu_6306_p1 = $unsigned(sext_ln142_34_fu_6302_p1);

assign zext_ln142_202_fu_6321_p1 = xor_ln899_103_fu_6315_p2;

assign zext_ln142_203_fu_6329_p1 = $unsigned(sext_ln142_35_fu_6325_p1);

assign zext_ln142_204_fu_6344_p1 = xor_ln899_104_fu_6338_p2;

assign zext_ln142_205_fu_6352_p1 = $unsigned(sext_ln142_36_fu_6348_p1);

assign zext_ln142_206_fu_6367_p1 = xor_ln899_105_fu_6361_p2;

assign zext_ln142_207_fu_6375_p1 = $unsigned(sext_ln142_37_fu_6371_p1);

assign zext_ln142_208_fu_6390_p1 = xor_ln899_106_fu_6384_p2;

assign zext_ln142_209_fu_6398_p1 = $unsigned(sext_ln142_38_fu_6394_p1);

assign zext_ln142_20_fu_4414_p1 = $unsigned(sext_ln142_1_fu_4410_p1);

assign zext_ln142_210_fu_6413_p1 = xor_ln899_107_fu_6407_p2;

assign zext_ln142_211_fu_6421_p1 = $unsigned(sext_ln142_39_fu_6417_p1);

assign zext_ln142_212_fu_6436_p1 = xor_ln899_108_fu_6430_p2;

assign zext_ln142_213_fu_6444_p1 = $unsigned(sext_ln142_40_fu_6440_p1);

assign zext_ln142_214_fu_6459_p1 = xor_ln899_109_fu_6453_p2;

assign zext_ln142_215_fu_6467_p1 = $unsigned(sext_ln142_41_fu_6463_p1);

assign zext_ln142_216_fu_6482_p1 = xor_ln899_110_fu_6476_p2;

assign zext_ln142_217_fu_6490_p1 = $unsigned(sext_ln142_42_fu_6486_p1);

assign zext_ln142_218_fu_6505_p1 = xor_ln899_111_fu_6499_p2;

assign zext_ln142_219_fu_6513_p1 = $unsigned(sext_ln142_43_fu_6509_p1);

assign zext_ln142_21_fu_4429_p1 = xor_ln899_11_fu_4423_p2;

assign zext_ln142_220_fu_6528_p1 = xor_ln899_112_fu_6522_p2;

assign zext_ln142_221_fu_6536_p1 = $unsigned(sext_ln142_44_fu_6532_p1);

assign zext_ln142_222_fu_6551_p1 = xor_ln899_113_fu_6545_p2;

assign zext_ln142_223_fu_6559_p1 = $unsigned(sext_ln142_45_fu_6555_p1);

assign zext_ln142_224_fu_6574_p1 = xor_ln899_114_fu_6568_p2;

assign zext_ln142_225_fu_6582_p1 = $unsigned(sext_ln142_46_fu_6578_p1);

assign zext_ln142_226_fu_6597_p1 = xor_ln899_115_fu_6591_p2;

assign zext_ln142_227_fu_6605_p1 = $unsigned(sext_ln142_47_fu_6601_p1);

assign zext_ln142_228_fu_6620_p1 = xor_ln899_116_fu_6614_p2;

assign zext_ln142_229_fu_6628_p1 = $unsigned(sext_ln142_48_fu_6624_p1);

assign zext_ln142_22_fu_4437_p1 = $unsigned(sext_ln142_2_fu_4433_p1);

assign zext_ln142_230_fu_6643_p1 = xor_ln899_117_fu_6637_p2;

assign zext_ln142_231_fu_6651_p1 = $unsigned(sext_ln142_49_fu_6647_p1);

assign zext_ln142_232_fu_6666_p1 = xor_ln899_118_fu_6660_p2;

assign zext_ln142_233_fu_6674_p1 = $unsigned(sext_ln142_50_fu_6670_p1);

assign zext_ln142_234_fu_6689_p1 = xor_ln899_119_fu_6683_p2;

assign zext_ln142_235_fu_6697_p1 = $unsigned(sext_ln142_51_fu_6693_p1);

assign zext_ln142_236_fu_6712_p1 = xor_ln899_120_fu_6706_p2;

assign zext_ln142_237_fu_6720_p1 = $unsigned(sext_ln142_52_fu_6716_p1);

assign zext_ln142_238_fu_6735_p1 = xor_ln899_121_fu_6729_p2;

assign zext_ln142_239_fu_6743_p1 = $unsigned(sext_ln142_53_fu_6739_p1);

assign zext_ln142_23_fu_4452_p1 = xor_ln899_12_fu_4446_p2;

assign zext_ln142_240_fu_6758_p1 = xor_ln899_122_fu_6752_p2;

assign zext_ln142_241_fu_6766_p1 = $unsigned(sext_ln142_54_fu_6762_p1);

assign zext_ln142_242_fu_6781_p1 = xor_ln899_123_fu_6775_p2;

assign zext_ln142_243_fu_6789_p1 = $unsigned(sext_ln142_55_fu_6785_p1);

assign zext_ln142_244_fu_6804_p1 = xor_ln899_124_fu_6798_p2;

assign zext_ln142_245_fu_6812_p1 = $unsigned(sext_ln142_56_fu_6808_p1);

assign zext_ln142_246_fu_6827_p1 = xor_ln899_125_fu_6821_p2;

assign zext_ln142_247_fu_6850_p1 = xor_ln899_126_fu_6844_p2;

assign zext_ln142_248_fu_6865_p1 = xor_ln899_127_fu_6859_p2;

assign zext_ln142_249_fu_6880_p1 = xor_ln899_128_fu_6874_p2;

assign zext_ln142_24_fu_4460_p1 = $unsigned(sext_ln142_3_fu_4456_p1);

assign zext_ln142_250_fu_6895_p1 = xor_ln899_129_fu_6889_p2;

assign zext_ln142_251_fu_6910_p1 = xor_ln899_130_fu_6904_p2;

assign zext_ln142_252_fu_6925_p1 = xor_ln899_131_fu_6919_p2;

assign zext_ln142_253_fu_6940_p1 = xor_ln899_132_fu_6934_p2;

assign zext_ln142_254_fu_6955_p1 = xor_ln899_133_fu_6949_p2;

assign zext_ln142_255_fu_6970_p1 = xor_ln899_134_fu_6964_p2;

assign zext_ln142_256_fu_6985_p1 = xor_ln899_135_fu_6979_p2;

assign zext_ln142_257_fu_7000_p1 = xor_ln899_136_fu_6994_p2;

assign zext_ln142_258_fu_7015_p1 = xor_ln899_137_fu_7009_p2;

assign zext_ln142_259_fu_7030_p1 = xor_ln899_138_fu_7024_p2;

assign zext_ln142_25_fu_4475_p1 = xor_ln899_13_fu_4469_p2;

assign zext_ln142_260_fu_7045_p1 = xor_ln899_139_fu_7039_p2;

assign zext_ln142_261_fu_7060_p1 = xor_ln899_140_fu_7054_p2;

assign zext_ln142_262_fu_7075_p1 = xor_ln899_141_fu_7069_p2;

assign zext_ln142_263_fu_7090_p1 = xor_ln899_142_fu_7084_p2;

assign zext_ln142_264_fu_7105_p1 = xor_ln899_143_fu_7099_p2;

assign zext_ln142_265_fu_7120_p1 = xor_ln899_144_fu_7114_p2;

assign zext_ln142_266_fu_7135_p1 = xor_ln899_145_fu_7129_p2;

assign zext_ln142_267_fu_7150_p1 = xor_ln899_146_fu_7144_p2;

assign zext_ln142_268_fu_7165_p1 = xor_ln899_147_fu_7159_p2;

assign zext_ln142_269_fu_7180_p1 = xor_ln899_148_fu_7174_p2;

assign zext_ln142_26_fu_4498_p1 = xor_ln899_14_fu_4492_p2;

assign zext_ln142_270_fu_7195_p1 = xor_ln899_149_fu_7189_p2;

assign zext_ln142_271_fu_7210_p1 = xor_ln899_150_fu_7204_p2;

assign zext_ln142_272_fu_7225_p1 = xor_ln899_151_fu_7219_p2;

assign zext_ln142_273_fu_7240_p1 = xor_ln899_152_fu_7234_p2;

assign zext_ln142_274_fu_7255_p1 = xor_ln899_153_fu_7249_p2;

assign zext_ln142_275_fu_7270_p1 = xor_ln899_154_fu_7264_p2;

assign zext_ln142_276_fu_7285_p1 = xor_ln899_155_fu_7279_p2;

assign zext_ln142_277_fu_7300_p1 = xor_ln899_156_fu_7294_p2;

assign zext_ln142_278_fu_7315_p1 = xor_ln899_157_fu_7309_p2;

assign zext_ln142_279_fu_7330_p1 = xor_ln899_158_fu_7324_p2;

assign zext_ln142_27_fu_4502_p1 = threshs_m_thresholds_197_q0;

assign zext_ln142_280_fu_7345_p1 = xor_ln899_159_fu_7339_p2;

assign zext_ln142_281_fu_7360_p1 = xor_ln899_160_fu_7354_p2;

assign zext_ln142_282_fu_7375_p1 = xor_ln899_161_fu_7369_p2;

assign zext_ln142_283_fu_7390_p1 = xor_ln899_162_fu_7384_p2;

assign zext_ln142_284_fu_7405_p1 = xor_ln899_163_fu_7399_p2;

assign zext_ln142_285_fu_7420_p1 = xor_ln899_164_fu_7414_p2;

assign zext_ln142_286_fu_7435_p1 = xor_ln899_165_fu_7429_p2;

assign zext_ln142_287_fu_7450_p1 = xor_ln899_166_fu_7444_p2;

assign zext_ln142_288_fu_7465_p1 = xor_ln899_167_fu_7459_p2;

assign zext_ln142_289_fu_7480_p1 = xor_ln899_168_fu_7474_p2;

assign zext_ln142_28_fu_4517_p1 = xor_ln899_15_fu_4511_p2;

assign zext_ln142_290_fu_7495_p1 = xor_ln899_169_fu_7489_p2;

assign zext_ln142_291_fu_7510_p1 = xor_ln899_170_fu_7504_p2;

assign zext_ln142_292_fu_7525_p1 = xor_ln899_171_fu_7519_p2;

assign zext_ln142_293_fu_7540_p1 = xor_ln899_172_fu_7534_p2;

assign zext_ln142_294_fu_7555_p1 = xor_ln899_173_fu_7549_p2;

assign zext_ln142_295_fu_7570_p1 = xor_ln899_174_fu_7564_p2;

assign zext_ln142_296_fu_7585_p1 = xor_ln899_175_fu_7579_p2;

assign zext_ln142_297_fu_7600_p1 = xor_ln899_176_fu_7594_p2;

assign zext_ln142_298_fu_7615_p1 = xor_ln899_177_fu_7609_p2;

assign zext_ln142_299_fu_7630_p1 = xor_ln899_178_fu_7624_p2;

assign zext_ln142_29_fu_4521_p1 = threshs_m_thresholds_186_q0;

assign zext_ln142_2_fu_4228_p1 = threshs_m_thresholds_253_q0;

assign zext_ln142_300_fu_7645_p1 = xor_ln899_179_fu_7639_p2;

assign zext_ln142_301_fu_7660_p1 = xor_ln899_180_fu_7654_p2;

assign zext_ln142_302_fu_7675_p1 = xor_ln899_181_fu_7669_p2;

assign zext_ln142_303_fu_7690_p1 = xor_ln899_182_fu_7684_p2;

assign zext_ln142_304_fu_7705_p1 = xor_ln899_183_fu_7699_p2;

assign zext_ln142_305_fu_7720_p1 = xor_ln899_184_fu_7714_p2;

assign zext_ln142_306_fu_7735_p1 = xor_ln899_185_fu_7729_p2;

assign zext_ln142_307_fu_7750_p1 = xor_ln899_186_fu_7744_p2;

assign zext_ln142_308_fu_7765_p1 = xor_ln899_187_fu_7759_p2;

assign zext_ln142_309_fu_7780_p1 = xor_ln899_188_fu_7774_p2;

assign zext_ln142_30_fu_4536_p1 = xor_ln899_16_fu_4530_p2;

assign zext_ln142_310_fu_7795_p1 = xor_ln899_189_fu_7789_p2;

assign zext_ln142_311_fu_7810_p1 = xor_ln899_190_fu_7804_p2;

assign zext_ln142_312_fu_7825_p1 = xor_ln899_191_fu_7819_p2;

assign zext_ln142_313_fu_7844_p1 = xor_ln899_192_fu_7838_p2;

assign zext_ln142_314_fu_7863_p1 = xor_ln899_193_fu_7857_p2;

assign zext_ln142_315_fu_7882_p1 = xor_ln899_194_fu_7876_p2;

assign zext_ln142_316_fu_7901_p1 = xor_ln899_195_fu_7895_p2;

assign zext_ln142_317_fu_7920_p1 = xor_ln899_196_fu_7914_p2;

assign zext_ln142_318_fu_7939_p1 = xor_ln899_197_fu_7933_p2;

assign zext_ln142_319_fu_7958_p1 = xor_ln899_198_fu_7952_p2;

assign zext_ln142_31_fu_4540_p1 = threshs_m_thresholds_175_q0;

assign zext_ln142_320_fu_7977_p1 = xor_ln899_199_fu_7971_p2;

assign zext_ln142_321_fu_7996_p1 = xor_ln899_200_fu_7990_p2;

assign zext_ln142_322_fu_8015_p1 = xor_ln899_201_fu_8009_p2;

assign zext_ln142_323_fu_8034_p1 = xor_ln899_202_fu_8028_p2;

assign zext_ln142_324_fu_8053_p1 = xor_ln899_203_fu_8047_p2;

assign zext_ln142_325_fu_8072_p1 = xor_ln899_204_fu_8066_p2;

assign zext_ln142_326_fu_8091_p1 = xor_ln899_205_fu_8085_p2;

assign zext_ln142_327_fu_8110_p1 = xor_ln899_206_fu_8104_p2;

assign zext_ln142_328_fu_8129_p1 = xor_ln899_207_fu_8123_p2;

assign zext_ln142_329_fu_8148_p1 = xor_ln899_208_fu_8142_p2;

assign zext_ln142_32_fu_4555_p1 = xor_ln899_17_fu_4549_p2;

assign zext_ln142_330_fu_8167_p1 = xor_ln899_209_fu_8161_p2;

assign zext_ln142_331_fu_8186_p1 = xor_ln899_210_fu_8180_p2;

assign zext_ln142_332_fu_8205_p1 = xor_ln899_211_fu_8199_p2;

assign zext_ln142_333_fu_8224_p1 = xor_ln899_212_fu_8218_p2;

assign zext_ln142_334_fu_8243_p1 = xor_ln899_213_fu_8237_p2;

assign zext_ln142_335_fu_8262_p1 = xor_ln899_214_fu_8256_p2;

assign zext_ln142_336_fu_8281_p1 = xor_ln899_215_fu_8275_p2;

assign zext_ln142_337_fu_8300_p1 = xor_ln899_216_fu_8294_p2;

assign zext_ln142_338_fu_8319_p1 = xor_ln899_217_fu_8313_p2;

assign zext_ln142_339_fu_8338_p1 = xor_ln899_218_fu_8332_p2;

assign zext_ln142_33_fu_4559_p1 = threshs_m_thresholds_164_q0;

assign zext_ln142_340_fu_8357_p1 = xor_ln899_219_fu_8351_p2;

assign zext_ln142_341_fu_8376_p1 = xor_ln899_220_fu_8370_p2;

assign zext_ln142_342_fu_8395_p1 = xor_ln899_221_fu_8389_p2;

assign zext_ln142_343_fu_8414_p1 = xor_ln899_222_fu_8408_p2;

assign zext_ln142_344_fu_8433_p1 = xor_ln899_223_fu_8427_p2;

assign zext_ln142_345_fu_8452_p1 = xor_ln899_224_fu_8446_p2;

assign zext_ln142_346_fu_8471_p1 = xor_ln899_225_fu_8465_p2;

assign zext_ln142_347_fu_8490_p1 = xor_ln899_226_fu_8484_p2;

assign zext_ln142_348_fu_8509_p1 = xor_ln899_227_fu_8503_p2;

assign zext_ln142_349_fu_8528_p1 = xor_ln899_228_fu_8522_p2;

assign zext_ln142_34_fu_4574_p1 = xor_ln899_18_fu_4568_p2;

assign zext_ln142_350_fu_8547_p1 = xor_ln899_229_fu_8541_p2;

assign zext_ln142_351_fu_8566_p1 = xor_ln899_230_fu_8560_p2;

assign zext_ln142_352_fu_8585_p1 = xor_ln899_231_fu_8579_p2;

assign zext_ln142_353_fu_8604_p1 = xor_ln899_232_fu_8598_p2;

assign zext_ln142_354_fu_8623_p1 = xor_ln899_233_fu_8617_p2;

assign zext_ln142_355_fu_8642_p1 = xor_ln899_234_fu_8636_p2;

assign zext_ln142_356_fu_8661_p1 = xor_ln899_235_fu_8655_p2;

assign zext_ln142_357_fu_8680_p1 = xor_ln899_236_fu_8674_p2;

assign zext_ln142_358_fu_8699_p1 = xor_ln899_237_fu_8693_p2;

assign zext_ln142_359_fu_8718_p1 = xor_ln899_238_fu_8712_p2;

assign zext_ln142_35_fu_4578_p1 = threshs_m_thresholds_153_q0;

assign zext_ln142_360_fu_8737_p1 = xor_ln899_239_fu_8731_p2;

assign zext_ln142_361_fu_8756_p1 = xor_ln899_240_fu_8750_p2;

assign zext_ln142_362_fu_8775_p1 = xor_ln899_241_fu_8769_p2;

assign zext_ln142_363_fu_8794_p1 = xor_ln899_242_fu_8788_p2;

assign zext_ln142_364_fu_8813_p1 = xor_ln899_243_fu_8807_p2;

assign zext_ln142_365_fu_8832_p1 = xor_ln899_244_fu_8826_p2;

assign zext_ln142_366_fu_8851_p1 = xor_ln899_245_fu_8845_p2;

assign zext_ln142_367_fu_8870_p1 = xor_ln899_246_fu_8864_p2;

assign zext_ln142_368_fu_8889_p1 = xor_ln899_247_fu_8883_p2;

assign zext_ln142_369_fu_8908_p1 = xor_ln899_248_fu_8902_p2;

assign zext_ln142_36_fu_4593_p1 = xor_ln899_19_fu_4587_p2;

assign zext_ln142_370_fu_8927_p1 = xor_ln899_249_fu_8921_p2;

assign zext_ln142_371_fu_8946_p1 = xor_ln899_250_fu_8940_p2;

assign zext_ln142_372_fu_8965_p1 = xor_ln899_251_fu_8959_p2;

assign zext_ln142_373_fu_8984_p1 = xor_ln899_252_fu_8978_p2;

assign zext_ln142_374_fu_9003_p1 = xor_ln899_253_fu_8997_p2;

assign zext_ln142_37_fu_4597_p1 = threshs_m_thresholds_141_q0;

assign zext_ln142_38_fu_4612_p1 = xor_ln899_20_fu_4606_p2;

assign zext_ln142_39_fu_4616_p1 = threshs_m_thresholds_130_q0;

assign zext_ln142_3_fu_10682_p1 = xor_ln899_1_fu_10677_p2;

assign zext_ln142_40_fu_4631_p1 = xor_ln899_21_fu_4625_p2;

assign zext_ln142_41_fu_4635_p1 = threshs_m_thresholds_119_q0;

assign zext_ln142_42_fu_4650_p1 = xor_ln899_22_fu_4644_p2;

assign zext_ln142_43_fu_4658_p1 = $unsigned(sext_ln142_4_fu_4654_p1);

assign zext_ln142_44_fu_4673_p1 = xor_ln899_23_fu_4667_p2;

assign zext_ln142_45_fu_4681_p1 = $unsigned(sext_ln142_5_fu_4677_p1);

assign zext_ln142_46_fu_4696_p1 = xor_ln899_24_fu_4690_p2;

assign zext_ln142_47_fu_4704_p1 = $unsigned(sext_ln142_6_fu_4700_p1);

assign zext_ln142_48_fu_4719_p1 = xor_ln899_25_fu_4713_p2;

assign zext_ln142_49_fu_4727_p1 = $unsigned(sext_ln142_7_fu_4723_p1);

assign zext_ln142_4_fu_10691_p1 = xor_ln899_2_fu_10686_p2;

assign zext_ln142_50_fu_4742_p1 = xor_ln899_26_fu_4736_p2;

assign zext_ln142_51_fu_4750_p1 = $unsigned(sext_ln142_8_fu_4746_p1);

assign zext_ln142_52_fu_4765_p1 = xor_ln899_27_fu_4759_p2;

assign zext_ln142_53_fu_4773_p1 = $unsigned(sext_ln142_9_fu_4769_p1);

assign zext_ln142_54_fu_4788_p1 = xor_ln899_28_fu_4782_p2;

assign zext_ln142_55_fu_4796_p1 = $unsigned(sext_ln142_10_fu_4792_p1);

assign zext_ln142_56_fu_4811_p1 = xor_ln899_29_fu_4805_p2;

assign zext_ln142_57_fu_4834_p1 = xor_ln899_30_fu_4828_p2;

assign zext_ln142_58_fu_4838_p1 = threshs_m_thresholds_74_q0;

assign zext_ln142_59_fu_4853_p1 = xor_ln899_31_fu_4847_p2;

assign zext_ln142_5_fu_4250_p1 = threshs_m_thresholds_76_q0;

assign zext_ln142_60_fu_4857_p1 = threshs_m_thresholds_73_q0;

assign zext_ln142_61_fu_4872_p1 = xor_ln899_32_fu_4866_p2;

assign zext_ln142_62_fu_4876_p1 = threshs_m_thresholds_72_q0;

assign zext_ln142_63_fu_4891_p1 = xor_ln899_33_fu_4885_p2;

assign zext_ln142_64_fu_4895_p1 = threshs_m_thresholds_71_q0;

assign zext_ln142_65_fu_4910_p1 = xor_ln899_34_fu_4904_p2;

assign zext_ln142_66_fu_4914_p1 = threshs_m_thresholds_70_q0;

assign zext_ln142_67_fu_4929_p1 = xor_ln899_35_fu_4923_p2;

assign zext_ln142_68_fu_4933_p1 = threshs_m_thresholds_69_q0;

assign zext_ln142_69_fu_4948_p1 = xor_ln899_36_fu_4942_p2;

assign zext_ln142_6_fu_4265_p1 = xor_ln899_3_fu_4259_p2;

assign zext_ln142_70_fu_4952_p1 = threshs_m_thresholds_68_q0;

assign zext_ln142_71_fu_4967_p1 = xor_ln899_37_fu_4961_p2;

assign zext_ln142_72_fu_4971_p1 = threshs_m_thresholds_67_q0;

assign zext_ln142_73_fu_4986_p1 = xor_ln899_38_fu_4980_p2;

assign zext_ln142_74_fu_4990_p1 = threshs_m_thresholds_66_q0;

assign zext_ln142_75_fu_5005_p1 = xor_ln899_39_fu_4999_p2;

assign zext_ln142_76_fu_5009_p1 = threshs_m_thresholds_64_q0;

assign zext_ln142_77_fu_5024_p1 = xor_ln899_40_fu_5018_p2;

assign zext_ln142_78_fu_5028_p1 = threshs_m_thresholds_63_q0;

assign zext_ln142_79_fu_5043_p1 = xor_ln899_41_fu_5037_p2;

assign zext_ln142_7_fu_4269_p1 = threshs_m_thresholds_65_q0;

assign zext_ln142_80_fu_5047_p1 = threshs_m_thresholds_62_q0;

assign zext_ln142_81_fu_5062_p1 = xor_ln899_42_fu_5056_p2;

assign zext_ln142_82_fu_5066_p1 = threshs_m_thresholds_61_q0;

assign zext_ln142_83_fu_5081_p1 = xor_ln899_43_fu_5075_p2;

assign zext_ln142_84_fu_5085_p1 = threshs_m_thresholds_60_q0;

assign zext_ln142_85_fu_5100_p1 = xor_ln899_44_fu_5094_p2;

assign zext_ln142_86_fu_5104_p1 = threshs_m_thresholds_59_q0;

assign zext_ln142_87_fu_5119_p1 = xor_ln899_45_fu_5113_p2;

assign zext_ln142_88_fu_5123_p1 = threshs_m_thresholds_58_q0;

assign zext_ln142_89_fu_5138_p1 = xor_ln899_46_fu_5132_p2;

assign zext_ln142_8_fu_4284_p1 = xor_ln899_4_fu_4278_p2;

assign zext_ln142_90_fu_5146_p1 = $unsigned(sext_ln142_11_fu_5142_p1);

assign zext_ln142_91_fu_5161_p1 = xor_ln899_47_fu_5155_p2;

assign zext_ln142_92_fu_5169_p1 = $unsigned(sext_ln142_12_fu_5165_p1);

assign zext_ln142_93_fu_5184_p1 = xor_ln899_48_fu_5178_p2;

assign zext_ln142_94_fu_5192_p1 = $unsigned(sext_ln142_13_fu_5188_p1);

assign zext_ln142_95_fu_5207_p1 = xor_ln899_49_fu_5201_p2;

assign zext_ln142_96_fu_5215_p1 = $unsigned(sext_ln142_14_fu_5211_p1);

assign zext_ln142_97_fu_5230_p1 = xor_ln899_50_fu_5224_p2;

assign zext_ln142_98_fu_5238_p1 = $unsigned(sext_ln142_15_fu_5234_p1);

assign zext_ln142_99_fu_5253_p1 = xor_ln899_51_fu_5247_p2;

assign zext_ln142_9_fu_4292_p1 = $unsigned(sext_ln142_fu_4288_p1);

assign zext_ln142_fu_3940_p1 = nf_assign_reg_3906;

assign zext_ln700_100_fu_9718_p1 = add_ln700_104_fu_9712_p2;

assign zext_ln700_101_fu_10983_p1 = add_ln700_105_reg_13190;

assign zext_ln700_102_fu_10992_p1 = add_ln700_106_fu_10986_p2;

assign zext_ln700_103_fu_11002_p1 = add_ln700_107_fu_10996_p2;

assign zext_ln700_104_fu_9734_p1 = add_ln700_108_fu_9728_p2;

assign zext_ln700_105_fu_9744_p1 = add_ln700_109_fu_9738_p2;

assign zext_ln700_106_fu_11006_p1 = add_ln700_110_reg_13195;

assign zext_ln700_107_fu_9760_p1 = add_ln700_111_fu_9754_p2;

assign zext_ln700_108_fu_9770_p1 = add_ln700_112_fu_9764_p2;

assign zext_ln700_109_fu_11009_p1 = add_ln700_113_reg_13200;

assign zext_ln700_10_fu_10723_p1 = add_ln700_11_reg_13070;

assign zext_ln700_110_fu_11018_p1 = add_ln700_114_fu_11012_p2;

assign zext_ln700_111_fu_9786_p1 = add_ln700_115_fu_9780_p2;

assign zext_ln700_112_fu_9796_p1 = add_ln700_116_fu_9790_p2;

assign zext_ln700_113_fu_11022_p1 = add_ln700_117_reg_13205;

assign zext_ln700_114_fu_9812_p1 = add_ln700_118_fu_9806_p2;

assign zext_ln700_115_fu_9822_p1 = add_ln700_119_fu_9816_p2;

assign zext_ln700_116_fu_11025_p1 = add_ln700_120_reg_13210;

assign zext_ln700_117_fu_11034_p1 = add_ln700_121_fu_11028_p2;

assign zext_ln700_118_fu_11044_p1 = add_ln700_122_fu_11038_p2;

assign zext_ln700_119_fu_11054_p1 = add_ln700_123_fu_11048_p2;

assign zext_ln700_11_fu_10732_p1 = add_ln700_12_fu_10726_p2;

assign zext_ln700_120_fu_11469_p1 = add_ln700_124_reg_13390;

assign zext_ln700_121_fu_9838_p1 = add_ln700_126_fu_9832_p2;

assign zext_ln700_122_fu_9848_p1 = add_ln700_127_fu_9842_p2;

assign zext_ln700_123_fu_11064_p1 = add_ln700_128_reg_13215;

assign zext_ln700_124_fu_9864_p1 = add_ln700_129_fu_9858_p2;

assign zext_ln700_125_fu_9874_p1 = add_ln700_130_fu_9868_p2;

assign zext_ln700_126_fu_11067_p1 = add_ln700_131_reg_13220;

assign zext_ln700_127_fu_11076_p1 = add_ln700_132_fu_11070_p2;

assign zext_ln700_128_fu_9890_p1 = add_ln700_133_fu_9884_p2;

assign zext_ln700_129_fu_9900_p1 = add_ln700_134_fu_9894_p2;

assign zext_ln700_12_fu_9110_p1 = add_ln700_14_fu_9104_p2;

assign zext_ln700_130_fu_11080_p1 = add_ln700_135_reg_13225;

assign zext_ln700_131_fu_9916_p1 = add_ln700_136_fu_9910_p2;

assign zext_ln700_132_fu_9926_p1 = add_ln700_137_fu_9920_p2;

assign zext_ln700_133_fu_11083_p1 = add_ln700_138_reg_13230;

assign zext_ln700_134_fu_11092_p1 = add_ln700_139_fu_11086_p2;

assign zext_ln700_135_fu_11102_p1 = add_ln700_140_fu_11096_p2;

assign zext_ln700_136_fu_9942_p1 = add_ln700_141_fu_9936_p2;

assign zext_ln700_137_fu_9952_p1 = add_ln700_142_fu_9946_p2;

assign zext_ln700_138_fu_11106_p1 = add_ln700_143_reg_13235;

assign zext_ln700_139_fu_9968_p1 = add_ln700_144_fu_9962_p2;

assign zext_ln700_13_fu_9120_p1 = add_ln700_15_fu_9114_p2;

assign zext_ln700_140_fu_9978_p1 = add_ln700_145_fu_9972_p2;

assign zext_ln700_141_fu_11109_p1 = add_ln700_146_reg_13240;

assign zext_ln700_142_fu_11118_p1 = add_ln700_147_fu_11112_p2;

assign zext_ln700_143_fu_9994_p1 = add_ln700_148_fu_9988_p2;

assign zext_ln700_144_fu_10004_p1 = add_ln700_149_fu_9998_p2;

assign zext_ln700_145_fu_11122_p1 = add_ln700_150_reg_13245;

assign zext_ln700_146_fu_10020_p1 = add_ln700_151_fu_10014_p2;

assign zext_ln700_147_fu_10030_p1 = add_ln700_152_fu_10024_p2;

assign zext_ln700_148_fu_11125_p1 = add_ln700_153_reg_13250;

assign zext_ln700_149_fu_11134_p1 = add_ln700_154_fu_11128_p2;

assign zext_ln700_14_fu_10742_p1 = add_ln700_16_reg_13075;

assign zext_ln700_150_fu_11144_p1 = add_ln700_155_fu_11138_p2;

assign zext_ln700_151_fu_11154_p1 = add_ln700_156_fu_11148_p2;

assign zext_ln700_152_fu_10046_p1 = add_ln700_157_fu_10040_p2;

assign zext_ln700_153_fu_10056_p1 = add_ln700_158_fu_10050_p2;

assign zext_ln700_154_fu_11158_p1 = add_ln700_159_reg_13255;

assign zext_ln700_155_fu_10072_p1 = add_ln700_160_fu_10066_p2;

assign zext_ln700_156_fu_10082_p1 = add_ln700_161_fu_10076_p2;

assign zext_ln700_157_fu_11161_p1 = add_ln700_162_reg_13260;

assign zext_ln700_158_fu_11170_p1 = add_ln700_163_fu_11164_p2;

assign zext_ln700_159_fu_10098_p1 = add_ln700_164_fu_10092_p2;

assign zext_ln700_15_fu_9136_p1 = add_ln700_17_fu_9130_p2;

assign zext_ln700_160_fu_10108_p1 = add_ln700_165_fu_10102_p2;

assign zext_ln700_161_fu_11174_p1 = add_ln700_166_reg_13265;

assign zext_ln700_162_fu_10124_p1 = add_ln700_167_fu_10118_p2;

assign zext_ln700_163_fu_10134_p1 = add_ln700_168_fu_10128_p2;

assign zext_ln700_164_fu_11177_p1 = add_ln700_169_reg_13270;

assign zext_ln700_165_fu_11186_p1 = add_ln700_170_fu_11180_p2;

assign zext_ln700_166_fu_11196_p1 = add_ln700_171_fu_11190_p2;

assign zext_ln700_167_fu_10150_p1 = add_ln700_172_fu_10144_p2;

assign zext_ln700_168_fu_10160_p1 = add_ln700_173_fu_10154_p2;

assign zext_ln700_169_fu_11200_p1 = add_ln700_174_reg_13275;

assign zext_ln700_16_fu_9146_p1 = add_ln700_18_fu_9140_p2;

assign zext_ln700_170_fu_10176_p1 = add_ln700_175_fu_10170_p2;

assign zext_ln700_171_fu_10186_p1 = add_ln700_176_fu_10180_p2;

assign zext_ln700_172_fu_11203_p1 = add_ln700_177_reg_13280;

assign zext_ln700_173_fu_11212_p1 = add_ln700_178_fu_11206_p2;

assign zext_ln700_174_fu_10202_p1 = add_ln700_179_fu_10196_p2;

assign zext_ln700_175_fu_10212_p1 = add_ln700_180_fu_10206_p2;

assign zext_ln700_176_fu_11216_p1 = add_ln700_181_reg_13285;

assign zext_ln700_177_fu_10228_p1 = add_ln700_182_fu_10222_p2;

assign zext_ln700_178_fu_10238_p1 = add_ln700_183_fu_10232_p2;

assign zext_ln700_179_fu_11219_p1 = add_ln700_184_reg_13290;

assign zext_ln700_17_fu_10745_p1 = add_ln700_19_reg_13080;

assign zext_ln700_180_fu_11228_p1 = add_ln700_185_fu_11222_p2;

assign zext_ln700_181_fu_11238_p1 = add_ln700_186_fu_11232_p2;

assign zext_ln700_182_fu_11248_p1 = add_ln700_187_fu_11242_p2;

assign zext_ln700_183_fu_11478_p1 = add_ln700_188_reg_13395;

assign zext_ln700_184_fu_10254_p1 = add_ln700_189_fu_10248_p2;

assign zext_ln700_185_fu_10264_p1 = add_ln700_190_fu_10258_p2;

assign zext_ln700_186_fu_11258_p1 = add_ln700_191_reg_13295;

assign zext_ln700_187_fu_10280_p1 = add_ln700_192_fu_10274_p2;

assign zext_ln700_188_fu_10290_p1 = add_ln700_193_fu_10284_p2;

assign zext_ln700_189_fu_11261_p1 = add_ln700_194_reg_13300;

assign zext_ln700_18_fu_10754_p1 = add_ln700_20_fu_10748_p2;

assign zext_ln700_190_fu_11270_p1 = add_ln700_195_fu_11264_p2;

assign zext_ln700_191_fu_10306_p1 = add_ln700_196_fu_10300_p2;

assign zext_ln700_192_fu_10316_p1 = add_ln700_197_fu_10310_p2;

assign zext_ln700_193_fu_11274_p1 = add_ln700_198_reg_13305;

assign zext_ln700_194_fu_10332_p1 = add_ln700_199_fu_10326_p2;

assign zext_ln700_195_fu_10342_p1 = add_ln700_200_fu_10336_p2;

assign zext_ln700_196_fu_11277_p1 = add_ln700_201_reg_13310;

assign zext_ln700_197_fu_11286_p1 = add_ln700_202_fu_11280_p2;

assign zext_ln700_198_fu_11296_p1 = add_ln700_203_fu_11290_p2;

assign zext_ln700_199_fu_10358_p1 = add_ln700_204_fu_10352_p2;

assign zext_ln700_19_fu_9162_p1 = add_ln700_21_fu_9156_p2;

assign zext_ln700_1_fu_10701_p1 = add_ln700_fu_10695_p2;

assign zext_ln700_200_fu_10368_p1 = add_ln700_205_fu_10362_p2;

assign zext_ln700_201_fu_11300_p1 = add_ln700_206_reg_13315;

assign zext_ln700_202_fu_10384_p1 = add_ln700_207_fu_10378_p2;

assign zext_ln700_203_fu_10394_p1 = add_ln700_208_fu_10388_p2;

assign zext_ln700_204_fu_11303_p1 = add_ln700_209_reg_13320;

assign zext_ln700_205_fu_11312_p1 = add_ln700_210_fu_11306_p2;

assign zext_ln700_206_fu_10410_p1 = add_ln700_211_fu_10404_p2;

assign zext_ln700_207_fu_10420_p1 = add_ln700_212_fu_10414_p2;

assign zext_ln700_208_fu_11316_p1 = add_ln700_213_reg_13325;

assign zext_ln700_209_fu_10436_p1 = add_ln700_214_fu_10430_p2;

assign zext_ln700_20_fu_9172_p1 = add_ln700_22_fu_9166_p2;

assign zext_ln700_210_fu_10446_p1 = add_ln700_215_fu_10440_p2;

assign zext_ln700_211_fu_11319_p1 = add_ln700_216_reg_13330;

assign zext_ln700_212_fu_11328_p1 = add_ln700_217_fu_11322_p2;

assign zext_ln700_213_fu_11338_p1 = add_ln700_218_fu_11332_p2;

assign zext_ln700_214_fu_11348_p1 = add_ln700_219_fu_11342_p2;

assign zext_ln700_215_fu_10462_p1 = add_ln700_220_fu_10456_p2;

assign zext_ln700_216_fu_10472_p1 = add_ln700_221_fu_10466_p2;

assign zext_ln700_217_fu_11352_p1 = add_ln700_222_reg_13335;

assign zext_ln700_218_fu_10488_p1 = add_ln700_223_fu_10482_p2;

assign zext_ln700_219_fu_10498_p1 = add_ln700_224_fu_10492_p2;

assign zext_ln700_21_fu_10758_p1 = add_ln700_23_reg_13085;

assign zext_ln700_220_fu_11355_p1 = add_ln700_225_reg_13340;

assign zext_ln700_221_fu_11364_p1 = add_ln700_226_fu_11358_p2;

assign zext_ln700_222_fu_10514_p1 = add_ln700_227_fu_10508_p2;

assign zext_ln700_223_fu_10524_p1 = add_ln700_228_fu_10518_p2;

assign zext_ln700_224_fu_11368_p1 = add_ln700_229_reg_13345;

assign zext_ln700_225_fu_10540_p1 = add_ln700_230_fu_10534_p2;

assign zext_ln700_226_fu_10550_p1 = add_ln700_231_fu_10544_p2;

assign zext_ln700_227_fu_11371_p1 = add_ln700_232_reg_13350;

assign zext_ln700_228_fu_11380_p1 = add_ln700_233_fu_11374_p2;

assign zext_ln700_229_fu_11390_p1 = add_ln700_234_fu_11384_p2;

assign zext_ln700_22_fu_9188_p1 = add_ln700_24_fu_9182_p2;

assign zext_ln700_230_fu_10566_p1 = add_ln700_235_fu_10560_p2;

assign zext_ln700_231_fu_10576_p1 = add_ln700_236_fu_10570_p2;

assign zext_ln700_232_fu_11394_p1 = add_ln700_237_reg_13355;

assign zext_ln700_233_fu_10592_p1 = add_ln700_238_fu_10586_p2;

assign zext_ln700_234_fu_10602_p1 = add_ln700_239_fu_10596_p2;

assign zext_ln700_235_fu_11397_p1 = add_ln700_240_reg_13360;

assign zext_ln700_236_fu_11406_p1 = add_ln700_241_fu_11400_p2;

assign zext_ln700_237_fu_10618_p1 = add_ln700_242_fu_10612_p2;

assign zext_ln700_238_fu_10628_p1 = add_ln700_243_fu_10622_p2;

assign zext_ln700_239_fu_11410_p1 = add_ln700_244_reg_13365;

assign zext_ln700_23_fu_9198_p1 = add_ln700_25_fu_9192_p2;

assign zext_ln700_240_fu_10644_p1 = add_ln700_245_fu_10638_p2;

assign zext_ln700_241_fu_10654_p1 = add_ln700_246_fu_10648_p2;

assign zext_ln700_242_fu_11413_p1 = add_ln700_247_reg_13370;

assign zext_ln700_243_fu_11422_p1 = add_ln700_248_fu_11416_p2;

assign zext_ln700_244_fu_11432_p1 = add_ln700_249_fu_11426_p2;

assign zext_ln700_245_fu_11442_p1 = add_ln700_250_fu_11436_p2;

assign zext_ln700_246_fu_11481_p1 = add_ln700_251_reg_13400;

assign zext_ln700_24_fu_10761_p1 = add_ln700_26_reg_13090;

assign zext_ln700_25_fu_10770_p1 = add_ln700_27_fu_10764_p2;

assign zext_ln700_26_fu_11452_p1 = add_ln700_28_reg_13380;

assign zext_ln700_27_fu_9214_p1 = add_ln700_30_fu_9208_p2;

assign zext_ln700_28_fu_9224_p1 = add_ln700_31_fu_9218_p2;

assign zext_ln700_29_fu_10780_p1 = add_ln700_32_reg_13095;

assign zext_ln700_2_fu_9032_p1 = add_ln700_2_fu_9026_p2;

assign zext_ln700_30_fu_9240_p1 = add_ln700_33_fu_9234_p2;

assign zext_ln700_31_fu_9250_p1 = add_ln700_34_fu_9244_p2;

assign zext_ln700_32_fu_10783_p1 = add_ln700_35_reg_13100;

assign zext_ln700_33_fu_10792_p1 = add_ln700_36_fu_10786_p2;

assign zext_ln700_34_fu_9266_p1 = add_ln700_37_fu_9260_p2;

assign zext_ln700_35_fu_9276_p1 = add_ln700_38_fu_9270_p2;

assign zext_ln700_36_fu_10796_p1 = add_ln700_39_reg_13105;

assign zext_ln700_37_fu_9292_p1 = add_ln700_40_fu_9286_p2;

assign zext_ln700_38_fu_9302_p1 = add_ln700_41_fu_9296_p2;

assign zext_ln700_39_fu_10799_p1 = add_ln700_42_reg_13110;

assign zext_ln700_3_fu_9042_p1 = add_ln700_3_fu_9036_p2;

assign zext_ln700_40_fu_10808_p1 = add_ln700_43_fu_10802_p2;

assign zext_ln700_41_fu_10818_p1 = add_ln700_44_fu_10812_p2;

assign zext_ln700_42_fu_9318_p1 = add_ln700_45_fu_9312_p2;

assign zext_ln700_43_fu_9328_p1 = add_ln700_46_fu_9322_p2;

assign zext_ln700_44_fu_10822_p1 = add_ln700_47_reg_13115;

assign zext_ln700_45_fu_9344_p1 = add_ln700_48_fu_9338_p2;

assign zext_ln700_46_fu_9354_p1 = add_ln700_49_fu_9348_p2;

assign zext_ln700_47_fu_10825_p1 = add_ln700_50_reg_13120;

assign zext_ln700_48_fu_10834_p1 = add_ln700_51_fu_10828_p2;

assign zext_ln700_49_fu_9370_p1 = add_ln700_52_fu_9364_p2;

assign zext_ln700_4_fu_10711_p1 = add_ln700_4_reg_13060;

assign zext_ln700_50_fu_9380_p1 = add_ln700_53_fu_9374_p2;

assign zext_ln700_51_fu_10838_p1 = add_ln700_54_reg_13125;

assign zext_ln700_52_fu_9396_p1 = add_ln700_55_fu_9390_p2;

assign zext_ln700_53_fu_9406_p1 = add_ln700_56_fu_9400_p2;

assign zext_ln700_54_fu_10841_p1 = add_ln700_57_reg_13130;

assign zext_ln700_55_fu_10850_p1 = add_ln700_58_fu_10844_p2;

assign zext_ln700_56_fu_10860_p1 = add_ln700_59_fu_10854_p2;

assign zext_ln700_57_fu_11460_p1 = add_ln700_60_reg_13385;

assign zext_ln700_58_fu_9422_p1 = add_ln700_62_fu_9416_p2;

assign zext_ln700_59_fu_9432_p1 = add_ln700_63_fu_9426_p2;

assign zext_ln700_5_fu_9058_p1 = add_ln700_6_fu_9052_p2;

assign zext_ln700_60_fu_10870_p1 = add_ln700_64_reg_13135;

assign zext_ln700_61_fu_9448_p1 = add_ln700_65_fu_9442_p2;

assign zext_ln700_62_fu_9458_p1 = add_ln700_66_fu_9452_p2;

assign zext_ln700_63_fu_10873_p1 = add_ln700_67_reg_13140;

assign zext_ln700_64_fu_10882_p1 = add_ln700_68_fu_10876_p2;

assign zext_ln700_65_fu_9474_p1 = add_ln700_69_fu_9468_p2;

assign zext_ln700_66_fu_9484_p1 = add_ln700_70_fu_9478_p2;

assign zext_ln700_67_fu_10886_p1 = add_ln700_71_reg_13145;

assign zext_ln700_68_fu_9500_p1 = add_ln700_72_fu_9494_p2;

assign zext_ln700_69_fu_9510_p1 = add_ln700_73_fu_9504_p2;

assign zext_ln700_6_fu_9068_p1 = add_ln700_7_fu_9062_p2;

assign zext_ln700_70_fu_10889_p1 = add_ln700_74_reg_13150;

assign zext_ln700_71_fu_10898_p1 = add_ln700_75_fu_10892_p2;

assign zext_ln700_72_fu_10908_p1 = add_ln700_76_fu_10902_p2;

assign zext_ln700_73_fu_9526_p1 = add_ln700_77_fu_9520_p2;

assign zext_ln700_74_fu_9536_p1 = add_ln700_78_fu_9530_p2;

assign zext_ln700_75_fu_10912_p1 = add_ln700_79_reg_13155;

assign zext_ln700_76_fu_9552_p1 = add_ln700_80_fu_9546_p2;

assign zext_ln700_77_fu_9562_p1 = add_ln700_81_fu_9556_p2;

assign zext_ln700_78_fu_10915_p1 = add_ln700_82_reg_13160;

assign zext_ln700_79_fu_10924_p1 = add_ln700_83_fu_10918_p2;

assign zext_ln700_7_fu_10720_p1 = add_ln700_8_reg_13065;

assign zext_ln700_80_fu_9578_p1 = add_ln700_84_fu_9572_p2;

assign zext_ln700_81_fu_9588_p1 = add_ln700_85_fu_9582_p2;

assign zext_ln700_82_fu_10928_p1 = add_ln700_86_reg_13165;

assign zext_ln700_83_fu_9604_p1 = add_ln700_87_fu_9598_p2;

assign zext_ln700_84_fu_9614_p1 = add_ln700_88_fu_9608_p2;

assign zext_ln700_85_fu_10931_p1 = add_ln700_89_reg_13170;

assign zext_ln700_86_fu_10940_p1 = add_ln700_90_fu_10934_p2;

assign zext_ln700_87_fu_10950_p1 = add_ln700_91_fu_10944_p2;

assign zext_ln700_88_fu_10960_p1 = add_ln700_92_fu_10954_p2;

assign zext_ln700_89_fu_9630_p1 = add_ln700_93_fu_9624_p2;

assign zext_ln700_8_fu_9084_p1 = add_ln700_9_fu_9078_p2;

assign zext_ln700_90_fu_9640_p1 = add_ln700_94_fu_9634_p2;

assign zext_ln700_91_fu_10964_p1 = add_ln700_95_reg_13175;

assign zext_ln700_92_fu_9656_p1 = add_ln700_96_fu_9650_p2;

assign zext_ln700_93_fu_9666_p1 = add_ln700_97_fu_9660_p2;

assign zext_ln700_94_fu_10967_p1 = add_ln700_98_reg_13180;

assign zext_ln700_95_fu_10976_p1 = add_ln700_99_fu_10970_p2;

assign zext_ln700_96_fu_9682_p1 = add_ln700_100_fu_9676_p2;

assign zext_ln700_97_fu_9692_p1 = add_ln700_101_fu_9686_p2;

assign zext_ln700_98_fu_10980_p1 = add_ln700_102_reg_13185;

assign zext_ln700_99_fu_9708_p1 = add_ln700_103_fu_9702_p2;

assign zext_ln700_9_fu_9094_p1 = add_ln700_10_fu_9088_p2;

assign zext_ln700_fu_9022_p1 = xor_ln899_254_fu_9016_p2;

endmodule //Thresholding_Batch_0_Thresholding_Batch
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcocq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_Batcocq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcocq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_Batcocq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_Batcocq_rom Thresholding_Batch_1_Thresholding_Batcocq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actmb6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actmb6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actmb6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actmb6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actmb6_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actmb6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/584e/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccxx.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccxx_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccxx_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccxx(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccxx_rom Thresholding_Batch_0_Thresholding_Batccxx_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actvdy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actvdy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actvdy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actvdy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actvdy_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actvdy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/841a/StreamingFIFO_6.v


module StreamingFIFO_6(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [23:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [23:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(24)
)
StreamingFIFO_6_StreamingFIFO_6
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_ConvolutionInputGenerator_3_0/synth/finn_design_ConvolutionInputGenerator_3_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:ConvolutionInputGenerator_3:1.0
// IP Revision: 2101301315

(* X_CORE_INFO = "ConvolutionInputGenerator_3_ConvolutionInputGenerator_3,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_ConvolutionInputGenerator_3_0,ConvolutionInputGenerator_3_ConvolutionInputGenerator_3,{}" *)
(* CORE_GENERATION_INFO = "finn_design_ConvolutionInputGenerator_3_0,ConvolutionInputGenerator_3_ConvolutionInputGenerator_3,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=ConvolutionInputGenerator_3,x_ipVersion=1.0,x_ipCoreRevision=2101301315,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_ConvolutionInputGenerator_3_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 4, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [31 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 4, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [31 : 0] out_V_V_TDATA;

  ConvolutionInputGenerator_3_ConvolutionInputGenerator_3 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/584e/StreamingFIFO_17.v


module StreamingFIFO_17(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(16)
)
StreamingFIFO_17_StreamingFIFO_17
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_15_0/synth/finn_design_StreamingFIFO_15_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_15:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_15,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_15_0,StreamingFIFO_15,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_15_0,StreamingFIFO_15,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_15,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_15_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [31 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 4, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [31 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 4, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_15 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingDataWidthConverter_Batch_5_0/synth/finn_design_StreamingDataWidthConverter_Batch_5_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingDataWidthConverter_Batch_5:1.0
// IP Revision: 2101301321

(* X_CORE_INFO = "StreamingDataWidthConverter_Batch_5_StreamingDataWidthConverter_Batch_5,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingDataWidthConverter_Batch_5_0,StreamingDataWidthConverter_Batch_5_StreamingDataWidthConverter_Batch_5,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingDataWidthConverter_Batch_5_0,StreamingDataWidthConverter_Batch_5_StreamingDataWidthConverter_Batch_5,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingDataWidthConverter_Batch_5,x_ipVersion=1.0,x_ipCoreRevision=2101301321,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingDataWidthConverter_Batch_5_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;

  StreamingDataWidthConverter_Batch_5_StreamingDataWidthConverter_Batch_5 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_BatckbM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_BatckbM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_BatckbM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_BatckbM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_BatckbM_rom Thresholding_Batch_1_Thresholding_BatckbM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actg8j.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actg8j_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actg8j_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actg8j(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actg8j_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actg8j_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActDeQ.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActDeQ_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActDeQ_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActDeQ(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActDeQ_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActDeQ_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_17_0/synth/finn_design_StreamingFIFO_17_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_17:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_17,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_17_0,StreamingFIFO_17,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_17_0,StreamingFIFO_17,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_17,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_17_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_17 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_BatclbW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_BatclbW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_BatclbW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_BatclbW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_BatclbW_rom Thresholding_Batch_2_Thresholding_BatclbW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcfYi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 3;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcfYi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcfYi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd3;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcfYi_rom Thresholding_Batch_0_Thresholding_BatcfYi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_3_wstrm_0/synth/finn_design_StreamingFCLayer_Batch_3_wstrm_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:user:memstream:1.0
// IP Revision: 5

(* X_CORE_INFO = "memstream,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_3_wstrm_0,memstream,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_3_wstrm_0,memstream,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=user,x_ipName=memstream,x_ipVersion=1.0,x_ipCoreRevision=5,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED,CONFIG_EN=true,NSTREAMS=1,MEM_DEPTH=144,MEM_WIDTH=48,MEM_INIT=/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/,RAM_STYLE=auto,STRM0_WIDTH=48,STRM1_WIDTH=32,STRM2_WIDTH=32,STRM3_WIDTH=32,STRM4_WIDTH=32,STRM5_WIDTH=32,STRM0\
_DEPTH=144,STRM1_DEPTH=2304,STRM2_DEPTH=2304,STRM3_DEPTH=2304,STRM4_DEPTH=2304,STRM5_DEPTH=2304,STRM0_OFFSET=0,STRM1_OFFSET=2304,STRM2_OFFSET=4608,STRM3_OFFSET=6912,STRM4_OFFSET=9216,STRM5_OFFSET=11520,AXILITE_ADDR_WIDTH=11}" *)
(* IP_DEFINITION_SOURCE = "package_project" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_3_wstrm_0 (
  aclk,
  aresetn,
  awready,
  awvalid,
  awaddr,
  awprot,
  wready,
  wvalid,
  wdata,
  wstrb,
  bready,
  bvalid,
  bresp,
  arready,
  arvalid,
  araddr,
  arprot,
  rready,
  rvalid,
  rresp,
  rdata,
  m_axis_0_tready,
  m_axis_0_tvalid,
  m_axis_0_tdata
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aclk, ASSOCIATED_BUSIF m_axis_0:m_axis_1:m_axis_2:m_axis_3:m_axis_4:m_axis_5:s_axilite, ASSOCIATED_RESET aresetn, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 aclk CLK" *)
input wire aclk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aresetn, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 aresetn RST" *)
input wire aresetn;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWREADY" *)
output wire awready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWVALID" *)
input wire awvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWADDR" *)
input wire [10 : 0] awaddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWPROT" *)
input wire [2 : 0] awprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WREADY" *)
output wire wready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WVALID" *)
input wire wvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WDATA" *)
input wire [31 : 0] wdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WSTRB" *)
input wire [3 : 0] wstrb;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BREADY" *)
input wire bready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BVALID" *)
output wire bvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BRESP" *)
output wire [1 : 0] bresp;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARREADY" *)
output wire arready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARVALID" *)
input wire arvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARADDR" *)
input wire [10 : 0] araddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARPROT" *)
input wire [2 : 0] arprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RREADY" *)
input wire rready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RVALID" *)
output wire rvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RRESP" *)
output wire [1 : 0] rresp;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axilite, DATA_WIDTH 32, PROTOCOL AXI4LITE, FREQ_HZ 100000000.000000, ID_WIDTH 0, ADDR_WIDTH 11, AWUSER_WIDTH 0, ARUSER_WIDTH 0, WUSER_WIDTH 0, RUSER_WIDTH 0, BUSER_WIDTH 0, READ_WRITE_MODE READ_WRITE, HAS_BURST 0, HAS_LOCK 0, HAS_PROT 1, HAS_CACHE 0, HAS_QOS 0, HAS_REGION 0, HAS_WSTRB 1, HAS_BRESP 1, HAS_RRESP 1, SUPPORTS_NARROW_BURST 0, NUM_READ_OUTSTANDING 1, NUM_WRITE_OUTSTANDING 1, MAX_BURST_LENGTH 1, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, NUM_READ_THREADS 1, NUM_W\
RITE_THREADS 1, RUSER_BITS_PER_BYTE 0, WUSER_BITS_PER_BYTE 0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RDATA" *)
output wire [31 : 0] rdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TREADY" *)
input wire m_axis_0_tready;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TVALID" *)
output wire m_axis_0_tvalid;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME m_axis_0, TDATA_NUM_BYTES 6, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TDATA" *)
output wire [47 : 0] m_axis_0_tdata;

  memstream #(
    .CONFIG_EN(1'B1),
    .NSTREAMS(1),
    .MEM_DEPTH(144),
    .MEM_WIDTH(48),
    .MEM_INIT("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/"),
    .RAM_STYLE("auto"),
    .STRM0_WIDTH(48),
    .STRM1_WIDTH(32),
    .STRM2_WIDTH(32),
    .STRM3_WIDTH(32),
    .STRM4_WIDTH(32),
    .STRM5_WIDTH(32),
    .STRM0_DEPTH(144),
    .STRM1_DEPTH(2304),
    .STRM2_DEPTH(2304),
    .STRM3_DEPTH(2304),
    .STRM4_DEPTH(2304),
    .STRM5_DEPTH(2304),
    .STRM0_OFFSET(0),
    .STRM1_OFFSET(2304),
    .STRM2_OFFSET(4608),
    .STRM3_OFFSET(6912),
    .STRM4_OFFSET(9216),
    .STRM5_OFFSET(11520),
    .AXILITE_ADDR_WIDTH(11)
  ) inst (
    .aclk(aclk),
    .aresetn(aresetn),
    .awready(awready),
    .awvalid(awvalid),
    .awaddr(awaddr),
    .awprot(awprot),
    .wready(wready),
    .wvalid(wvalid),
    .wdata(wdata),
    .wstrb(wstrb),
    .bready(bready),
    .bvalid(bvalid),
    .bresp(bresp),
    .arready(arready),
    .arvalid(arvalid),
    .araddr(araddr),
    .arprot(arprot),
    .rready(rready),
    .rvalid(rvalid),
    .rresp(rresp),
    .rdata(rdata),
    .m_axis_0_afull(1'B0),
    .m_axis_0_tready(m_axis_0_tready),
    .m_axis_0_tvalid(m_axis_0_tvalid),
    .m_axis_0_tdata(m_axis_0_tdata),
    .m_axis_1_afull(1'B0),
    .m_axis_1_tready(1'B1),
    .m_axis_1_tvalid(),
    .m_axis_1_tdata(),
    .m_axis_2_afull(1'B0),
    .m_axis_2_tready(1'B1),
    .m_axis_2_tvalid(),
    .m_axis_2_tdata(),
    .m_axis_3_afull(1'B0),
    .m_axis_3_tready(1'B1),
    .m_axis_3_tvalid(),
    .m_axis_3_tdata(),
    .m_axis_4_afull(1'B0),
    .m_axis_4_tready(1'B1),
    .m_axis_4_tvalid(),
    .m_axis_4_tdata(),
    .m_axis_5_afull(1'B0),
    .m_axis_5_tready(1'B1),
    .m_axis_5_tvalid(),
    .m_axis_5_tdata()
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActPgM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActPgM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActPgM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActPgM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActPgM_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActPgM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccDy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccDy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccDy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccDy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccDy_rom Thresholding_Batch_0_Thresholding_BatccDy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccgu.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccgu_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccgu_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccgu(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccgu_rom Thresholding_Batch_0_Thresholding_Batccgu_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_13_0/synth/finn_design_StreamingFIFO_13_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_13:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_13,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_13_0,StreamingFIFO_13,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_13_0,StreamingFIFO_13,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_13,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_13_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [31 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 4, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [31 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 4, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_13 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbjl.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbjl_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbjl_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbjl(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbjl_rom Thresholding_Batch_0_Thresholding_Batcbjl_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/7fe4/hdl/verilog/StreamingDataWidthConverter_Batch_3_StreamingDataWidthCo_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingDataWidthConverter_Batch_3_StreamingDataWidthCo_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [15:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln402_fu_88_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln411_reg_154;
reg   [15:0] r_V_reg_61;
reg   [7:0] t_0_reg_72;
reg   [0:0] icmp_ln402_reg_135;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [7:0] t_fu_94_p2;
reg   [15:0] tmp_V_reg_144;
wire   [31:0] p_Result_s_fu_103_p3;
reg   [31:0] p_Result_s_reg_149;
wire   [0:0] icmp_ln411_fu_117_p2;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg   [15:0] ap_phi_mux_r_V_phi_fu_65_p4;
reg   [31:0] i_1_fu_44;
wire   [31:0] i_fu_111_p2;
reg    ap_block_pp0_stage0_01001;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_fu_117_p2 == 1'd0) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_1_fu_44 <= i_fu_111_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_fu_117_p2 == 1'd1) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        i_1_fu_44 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_reg_135 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        r_V_reg_61 <= tmp_V_reg_144;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        r_V_reg_61 <= 16'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        t_0_reg_72 <= t_fu_94_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        t_0_reg_72 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln402_reg_135 <= icmp_ln402_fu_88_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln411_reg_154 <= icmp_ln411_fu_117_p2;
        p_Result_s_reg_149 <= p_Result_s_fu_103_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_reg_144 <= in_V_V_TDATA;
    end
end

always @ (*) begin
    if ((icmp_ln402_fu_88_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln402_reg_135 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_r_V_phi_fu_65_p4 = tmp_V_reg_144;
    end else begin
        ap_phi_mux_r_V_phi_fu_65_p4 = r_V_reg_61;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln402_fu_88_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln411_reg_154 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_reg_154 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln402_fu_88_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln402_fu_88_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0));
end

always @ (*) begin
    ap_block_state3_io = ((icmp_ln411_reg_154 == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign i_fu_111_p2 = (i_1_fu_44 + 32'd1);

assign icmp_ln402_fu_88_p2 = ((t_0_reg_72 == 8'd128) ? 1'b1 : 1'b0);

assign icmp_ln411_fu_117_p2 = ((i_fu_111_p2 == 32'd2) ? 1'b1 : 1'b0);

assign out_V_V_TDATA = p_Result_s_reg_149;

assign p_Result_s_fu_103_p3 = {{in_V_V_TDATA}, {ap_phi_mux_r_V_phi_fu_65_p4}};

assign t_fu_94_p2 = (t_0_reg_72 + 8'd1);

endmodule //StreamingDataWidthConverter_Batch_3_StreamingDataWidthCo_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcRg6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcRg6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcRg6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcRg6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcRg6_rom Thresholding_Batch_0_Thresholding_BatcRg6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actibs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actibs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actibs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actibs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actibs_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actibs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_StreamingFCLayer_Batch_4.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingFCLayer_Batch_4_StreamingFCLayer_Batch_4,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.409000,HLS_SYN_LAT=8200,HLS_SYN_TPT=none,HLS_SYN_MEM=56,HLS_SYN_DSP=0,HLS_SYN_FF=2662,HLS_SYN_LUT=3233,HLS_VERSION=2020_1_1}" *)

module StreamingFCLayer_Batch_4_StreamingFCLayer_Batch_4 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        weights_V_V_TDATA,
        weights_V_V_TVALID,
        weights_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [31:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
input  [127:0] weights_V_V_TDATA;
input   weights_V_V_TVALID;
output   weights_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;
reg weights_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_Matrix_Vector_Activa_fu_140_ap_start;
wire    grp_Matrix_Vector_Activa_fu_140_ap_done;
wire    grp_Matrix_Vector_Activa_fu_140_ap_idle;
wire    grp_Matrix_Vector_Activa_fu_140_ap_ready;
wire    grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY;
wire   [15:0] grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA;
wire    grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID;
wire    grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY;
wire    grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY;
reg    grp_Matrix_Vector_Activa_fu_140_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [31:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    regslice_both_weights_V_V_U_apdone_blk;
wire   [127:0] weights_V_V_TDATA_int;
wire    weights_V_V_TVALID_int;
reg    weights_V_V_TREADY_int;
wire    regslice_both_weights_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_Matrix_Vector_Activa_fu_140_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingFCLayer_Batch_4_Matrix_Vector_Activa grp_Matrix_Vector_Activa_fu_140(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_Matrix_Vector_Activa_fu_140_ap_start),
    .ap_done(grp_Matrix_Vector_Activa_fu_140_ap_done),
    .ap_idle(grp_Matrix_Vector_Activa_fu_140_ap_idle),
    .ap_ready(grp_Matrix_Vector_Activa_fu_140_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY),
    .out_V_V_TDATA(grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA),
    .out_V_V_TVALID(grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID),
    .out_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY),
    .weight_V_V_TDATA(weights_V_V_TDATA_int),
    .weight_V_V_TVALID(weights_V_V_TVALID_int),
    .weight_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 32 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 128 ))
regslice_both_weights_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(weights_V_V_TDATA),
    .vld_in(weights_V_V_TVALID),
    .ack_in(regslice_both_weights_V_V_U_ack_in),
    .data_out(weights_V_V_TDATA_int),
    .vld_out(weights_V_V_TVALID_int),
    .ack_out(weights_V_V_TREADY_int),
    .apdone_blk(regslice_both_weights_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA),
    .vld_in(grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b1;
        end else if ((grp_Matrix_Vector_Activa_fu_140_ap_ready == 1'b1)) begin
            grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    if (((regslice_both_weights_V_V_U_ack_in == 1'b1) & (weights_V_V_TVALID == 1'b1))) begin
        weights_V_V_TREADY = 1'b1;
    end else begin
        weights_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        weights_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY;
    end else begin
        weights_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_Matrix_Vector_Activa_fu_140_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_Matrix_Vector_Activa_fu_140_ap_start = grp_Matrix_Vector_Activa_fu_140_ap_start_reg;

assign grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingFCLayer_Batch_4_StreamingFCLayer_Batch_4
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/1ba7/StreamingFIFO_12.v


module StreamingFIFO_12(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [31:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(32)
)
StreamingFIFO_12_StreamingFIFO_12
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_16_0/synth/finn_design_StreamingFIFO_16_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_16:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_16,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_16_0,StreamingFIFO_16,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_16_0,StreamingFIFO_16,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_16,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_16_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [7 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_16 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Act2iS.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Act2iS_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Act2iS_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Act2iS(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Act2iS_rom StreamingFCLayer_Batch_3_Matrix_Vector_Act2iS_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingDataWidthConverter_Batch_0_0/synth/finn_design_StreamingDataWidthConverter_Batch_0_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingDataWidthConverter_Batch_0:1.0
// IP Revision: 2101301323

(* X_CORE_INFO = "StreamingDataWidthConverter_Batch_0_StreamingDataWidthConverter_Batch_0,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingDataWidthConverter_Batch_0_0,StreamingDataWidthConverter_Batch_0_StreamingDataWidthConverter_Batch_0,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingDataWidthConverter_Batch_0_0,StreamingDataWidthConverter_Batch_0_StreamingDataWidthConverter_Batch_0,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingDataWidthConverter_Batch_0,x_ipVersion=1.0,x_ipCoreRevision=2101301323,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingDataWidthConverter_Batch_0_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [7 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 3, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [23 : 0] out_V_V_TDATA;

  StreamingDataWidthConverter_Batch_0_StreamingDataWidthConverter_Batch_0 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actyd2.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actyd2_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actyd2_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actyd2(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actyd2_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actyd2_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/6405/hdl/verilog/StreamingFCLayer_Batch_5_StreamingFCLayer_cud.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

(* use_dsp = "no" *) module StreamingFCLayer_Batch_5_StreamingFCLayer_cud_Mul_LUT_0(a, b, p);
input[4 - 1 : 0] a; 
input[4 - 1 : 0] b; 
output[8 - 1 : 0] p;

assign p = $signed(a) * $signed(b);
endmodule
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_5_StreamingFCLayer_cud(
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



StreamingFCLayer_Batch_5_StreamingFCLayer_cud_Mul_LUT_0 StreamingFCLayer_Batch_5_StreamingFCLayer_cud_Mul_LUT_0_U(
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdeE_x.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcdeE_x_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdeE_x_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcdeE_x(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcdeE_x_rom Thresholding_Batch_0_Thresholding_BatcdeE_x_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4c0f/hdl/verilog/StreamingDataWidthConverter_Batch_0_StreamingDataWidthCo_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingDataWidthConverter_Batch_0_StreamingDataWidthCo_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [7:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [23:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln402_fu_96_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln411_reg_175;
reg   [15:0] r_V_reg_69;
reg   [11:0] t_0_reg_80;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [11:0] t_fu_102_p2;
wire   [23:0] p_Result_s_fu_111_p3;
reg   [23:0] p_Result_s_reg_170;
wire   [0:0] icmp_ln411_fu_125_p2;
wire   [15:0] trunc_ln_fu_146_p3;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg   [31:0] i_1_fu_52;
wire   [31:0] i_fu_119_p2;
reg    ap_block_pp0_stage0_01001;
wire   [7:0] tmp_1_fu_136_p4;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_fu_125_p2 == 1'd0) & (icmp_ln402_fu_96_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_1_fu_52 <= i_fu_119_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_fu_125_p2 == 1'd1) & (icmp_ln402_fu_96_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        i_1_fu_52 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_96_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        r_V_reg_69 <= trunc_ln_fu_146_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        r_V_reg_69 <= 16'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_96_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        t_0_reg_80 <= t_fu_102_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        t_0_reg_80 <= 12'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_96_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln411_reg_175 <= icmp_ln411_fu_125_p2;
        p_Result_s_reg_170 <= p_Result_s_fu_111_p3;
    end
end

always @ (*) begin
    if ((icmp_ln402_fu_96_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln402_fu_96_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_96_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln411_reg_175 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_reg_175 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln402_fu_96_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln402_fu_96_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((icmp_ln402_fu_96_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((icmp_ln402_fu_96_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((icmp_ln402_fu_96_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = ((icmp_ln402_fu_96_p2 == 1'd0) & (in_V_V_TVALID == 1'b0));
end

always @ (*) begin
    ap_block_state3_io = ((icmp_ln411_reg_175 == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign i_fu_119_p2 = (i_1_fu_52 + 32'd1);

assign icmp_ln402_fu_96_p2 = ((t_0_reg_80 == 12'd3072) ? 1'b1 : 1'b0);

assign icmp_ln411_fu_125_p2 = ((i_fu_119_p2 == 32'd3) ? 1'b1 : 1'b0);

assign out_V_V_TDATA = p_Result_s_reg_170;

assign p_Result_s_fu_111_p3 = {{in_V_V_TDATA}, {r_V_reg_69}};

assign t_fu_102_p2 = (t_0_reg_80 + 12'd1);

assign tmp_1_fu_136_p4 = {{r_V_reg_69[15:8]}};

assign trunc_ln_fu_146_p3 = {{in_V_V_TDATA}, {tmp_1_fu_136_p4}};

endmodule //StreamingDataWidthConverter_Batch_0_StreamingDataWidthCo_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActEe0.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActEe0_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActEe0_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActEe0(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActEe0_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActEe0_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActfYi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActfYi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActfYi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActfYi_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActfYi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActxdS.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActxdS_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActxdS_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActxdS(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActxdS_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActxdS_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActWhU.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActWhU_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActWhU_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActWhU(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActWhU_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActWhU_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbnm.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbnm_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbnm_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbnm(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbnm_rom Thresholding_Batch_0_Thresholding_Batcbnm_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccjv.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccjv_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccjv_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccjv(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccjv_rom Thresholding_Batch_0_Thresholding_Batccjv_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actocq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actocq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actocq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actocq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actocq_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actocq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Act4jc.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Act4jc_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Act4jc_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Act4jc(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Act4jc_rom StreamingFCLayer_Batch_2_Matrix_Vector_Act4jc_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actocq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actocq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actocq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actocq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actocq_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actocq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActIfE.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActIfE_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActIfE_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActIfE(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActIfE_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActIfE_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/cd9c/hdl/verilog/StreamingFCLayer_Batch_0_StreamingFCLayer_bkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module StreamingFCLayer_Batch_0_StreamingFCLayer_bkb #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH       = 32,
    din5_WIDTH       = 32,
    din6_WIDTH       = 32,
    din7_WIDTH       = 32,
    din8_WIDTH       = 32,
    din9_WIDTH       = 32,
    din10_WIDTH       = 32,
    din11_WIDTH       = 32,
    din12_WIDTH       = 32,
    din13_WIDTH       = 32,
    din14_WIDTH       = 32,
    din15_WIDTH       = 32,
    din16_WIDTH       = 32,
    din17_WIDTH       = 32,
    din18_WIDTH       = 32,
    din19_WIDTH       = 32,
    din20_WIDTH       = 32,
    din21_WIDTH       = 32,
    din22_WIDTH       = 32,
    din23_WIDTH       = 32,
    din24_WIDTH       = 32,
    din25_WIDTH       = 32,
    din26_WIDTH       = 32,
    din27_WIDTH       = 32,
    din28_WIDTH       = 32,
    din29_WIDTH       = 32,
    din30_WIDTH       = 32,
    din31_WIDTH       = 32,
    din32_WIDTH       = 32,
    din33_WIDTH       = 32,
    din34_WIDTH       = 32,
    din35_WIDTH       = 32,
    din36_WIDTH       = 32,
    din37_WIDTH       = 32,
    din38_WIDTH       = 32,
    din39_WIDTH       = 32,
    din40_WIDTH       = 32,
    din41_WIDTH       = 32,
    din42_WIDTH       = 32,
    din43_WIDTH       = 32,
    din44_WIDTH       = 32,
    din45_WIDTH       = 32,
    din46_WIDTH       = 32,
    din47_WIDTH       = 32,
    din48_WIDTH       = 32,
    din49_WIDTH       = 32,
    din50_WIDTH       = 32,
    din51_WIDTH       = 32,
    din52_WIDTH       = 32,
    din53_WIDTH       = 32,
    din54_WIDTH       = 32,
    din55_WIDTH       = 32,
    din56_WIDTH       = 32,
    din57_WIDTH       = 32,
    din58_WIDTH       = 32,
    din59_WIDTH       = 32,
    din60_WIDTH       = 32,
    din61_WIDTH       = 32,
    din62_WIDTH       = 32,
    din63_WIDTH       = 32,
    din64_WIDTH       = 32,
    din65_WIDTH       = 32,
    din66_WIDTH       = 32,
    din67_WIDTH       = 32,
    din68_WIDTH       = 32,
    din69_WIDTH       = 32,
    din70_WIDTH       = 32,
    din71_WIDTH       = 32,
    din72_WIDTH       = 32,
    din73_WIDTH       = 32,
    din74_WIDTH       = 32,
    din75_WIDTH       = 32,
    din76_WIDTH       = 32,
    din77_WIDTH       = 32,
    din78_WIDTH       = 32,
    din79_WIDTH       = 32,
    din80_WIDTH       = 32,
    din81_WIDTH       = 32,
    din82_WIDTH       = 32,
    din83_WIDTH       = 32,
    din84_WIDTH       = 32,
    din85_WIDTH       = 32,
    din86_WIDTH       = 32,
    din87_WIDTH       = 32,
    din88_WIDTH       = 32,
    din89_WIDTH       = 32,
    din90_WIDTH       = 32,
    din91_WIDTH       = 32,
    din92_WIDTH       = 32,
    din93_WIDTH       = 32,
    din94_WIDTH       = 32,
    din95_WIDTH       = 32,
    din96_WIDTH       = 32,
    din97_WIDTH       = 32,
    din98_WIDTH       = 32,
    din99_WIDTH       = 32,
    din100_WIDTH       = 32,
    din101_WIDTH       = 32,
    din102_WIDTH       = 32,
    din103_WIDTH       = 32,
    din104_WIDTH       = 32,
    din105_WIDTH       = 32,
    din106_WIDTH       = 32,
    din107_WIDTH       = 32,
    din108_WIDTH       = 32,
    din109_WIDTH       = 32,
    din110_WIDTH       = 32,
    din111_WIDTH       = 32,
    din112_WIDTH       = 32,
    din113_WIDTH       = 32,
    din114_WIDTH       = 32,
    din115_WIDTH       = 32,
    din116_WIDTH       = 32,
    din117_WIDTH       = 32,
    din118_WIDTH       = 32,
    din119_WIDTH       = 32,
    din120_WIDTH       = 32,
    din121_WIDTH       = 32,
    din122_WIDTH       = 32,
    din123_WIDTH       = 32,
    din124_WIDTH       = 32,
    din125_WIDTH       = 32,
    din126_WIDTH       = 32,
    din127_WIDTH       = 32,
    din128_WIDTH       = 32,
    din129_WIDTH       = 32,
    din130_WIDTH       = 32,
    din131_WIDTH       = 32,
    din132_WIDTH       = 32,
    din133_WIDTH       = 32,
    din134_WIDTH       = 32,
    din135_WIDTH       = 32,
    din136_WIDTH       = 32,
    din137_WIDTH       = 32,
    din138_WIDTH       = 32,
    din139_WIDTH       = 32,
    din140_WIDTH       = 32,
    din141_WIDTH       = 32,
    din142_WIDTH       = 32,
    din143_WIDTH       = 32,
    din144_WIDTH       = 32,
    din145_WIDTH       = 32,
    din146_WIDTH       = 32,
    din147_WIDTH       = 32,
    din148_WIDTH       = 32,
    din149_WIDTH       = 32,
    din150_WIDTH       = 32,
    din151_WIDTH       = 32,
    din152_WIDTH       = 32,
    din153_WIDTH       = 32,
    din154_WIDTH       = 32,
    din155_WIDTH       = 32,
    din156_WIDTH       = 32,
    din157_WIDTH       = 32,
    din158_WIDTH       = 32,
    din159_WIDTH       = 32,
    din160_WIDTH       = 32,
    din161_WIDTH       = 32,
    din162_WIDTH       = 32,
    din163_WIDTH       = 32,
    din164_WIDTH       = 32,
    din165_WIDTH       = 32,
    din166_WIDTH       = 32,
    din167_WIDTH       = 32,
    din168_WIDTH       = 32,
    din169_WIDTH       = 32,
    din170_WIDTH       = 32,
    din171_WIDTH       = 32,
    din172_WIDTH       = 32,
    din173_WIDTH       = 32,
    din174_WIDTH       = 32,
    din175_WIDTH       = 32,
    din176_WIDTH       = 32,
    din177_WIDTH       = 32,
    din178_WIDTH       = 32,
    din179_WIDTH       = 32,
    din180_WIDTH       = 32,
    din181_WIDTH       = 32,
    din182_WIDTH       = 32,
    din183_WIDTH       = 32,
    din184_WIDTH       = 32,
    din185_WIDTH       = 32,
    din186_WIDTH       = 32,
    din187_WIDTH       = 32,
    din188_WIDTH       = 32,
    din189_WIDTH       = 32,
    din190_WIDTH       = 32,
    din191_WIDTH       = 32,
    din192_WIDTH       = 32,
    din193_WIDTH       = 32,
    din194_WIDTH       = 32,
    din195_WIDTH       = 32,
    din196_WIDTH       = 32,
    din197_WIDTH       = 32,
    din198_WIDTH       = 32,
    din199_WIDTH       = 32,
    din200_WIDTH       = 32,
    din201_WIDTH       = 32,
    din202_WIDTH       = 32,
    din203_WIDTH       = 32,
    din204_WIDTH       = 32,
    din205_WIDTH       = 32,
    din206_WIDTH       = 32,
    din207_WIDTH       = 32,
    din208_WIDTH       = 32,
    din209_WIDTH       = 32,
    din210_WIDTH       = 32,
    din211_WIDTH       = 32,
    din212_WIDTH       = 32,
    din213_WIDTH       = 32,
    din214_WIDTH       = 32,
    din215_WIDTH       = 32,
    din216_WIDTH       = 32,
    din217_WIDTH       = 32,
    din218_WIDTH       = 32,
    din219_WIDTH       = 32,
    din220_WIDTH       = 32,
    din221_WIDTH       = 32,
    din222_WIDTH       = 32,
    din223_WIDTH       = 32,
    din224_WIDTH       = 32,
    din225_WIDTH       = 32,
    din226_WIDTH       = 32,
    din227_WIDTH       = 32,
    din228_WIDTH       = 32,
    din229_WIDTH       = 32,
    din230_WIDTH       = 32,
    din231_WIDTH       = 32,
    din232_WIDTH       = 32,
    din233_WIDTH       = 32,
    din234_WIDTH       = 32,
    din235_WIDTH       = 32,
    din236_WIDTH       = 32,
    din237_WIDTH       = 32,
    din238_WIDTH       = 32,
    din239_WIDTH       = 32,
    din240_WIDTH       = 32,
    din241_WIDTH       = 32,
    din242_WIDTH       = 32,
    din243_WIDTH       = 32,
    din244_WIDTH       = 32,
    din245_WIDTH       = 32,
    din246_WIDTH       = 32,
    din247_WIDTH       = 32,
    din248_WIDTH       = 32,
    din249_WIDTH       = 32,
    din250_WIDTH       = 32,
    din251_WIDTH       = 32,
    din252_WIDTH       = 32,
    din253_WIDTH       = 32,
    din254_WIDTH       = 32,
    din255_WIDTH       = 32,
    din256_WIDTH       = 32,
    din257_WIDTH       = 32,
    din258_WIDTH       = 32,
    din259_WIDTH       = 32,
    din260_WIDTH       = 32,
    din261_WIDTH       = 32,
    din262_WIDTH       = 32,
    din263_WIDTH       = 32,
    din264_WIDTH       = 32,
    din265_WIDTH       = 32,
    din266_WIDTH       = 32,
    din267_WIDTH       = 32,
    din268_WIDTH       = 32,
    din269_WIDTH       = 32,
    din270_WIDTH       = 32,
    din271_WIDTH       = 32,
    din272_WIDTH       = 32,
    din273_WIDTH       = 32,
    din274_WIDTH       = 32,
    din275_WIDTH       = 32,
    din276_WIDTH       = 32,
    din277_WIDTH       = 32,
    din278_WIDTH       = 32,
    din279_WIDTH       = 32,
    din280_WIDTH       = 32,
    din281_WIDTH       = 32,
    din282_WIDTH       = 32,
    din283_WIDTH       = 32,
    din284_WIDTH       = 32,
    din285_WIDTH       = 32,
    din286_WIDTH       = 32,
    din287_WIDTH       = 32,
    din288_WIDTH       = 32,
    din289_WIDTH       = 32,
    din290_WIDTH       = 32,
    din291_WIDTH       = 32,
    din292_WIDTH       = 32,
    din293_WIDTH       = 32,
    din294_WIDTH       = 32,
    din295_WIDTH       = 32,
    din296_WIDTH       = 32,
    din297_WIDTH       = 32,
    din298_WIDTH       = 32,
    din299_WIDTH       = 32,
    din300_WIDTH       = 32,
    din301_WIDTH       = 32,
    din302_WIDTH       = 32,
    din303_WIDTH       = 32,
    din304_WIDTH       = 32,
    din305_WIDTH       = 32,
    din306_WIDTH       = 32,
    din307_WIDTH       = 32,
    din308_WIDTH       = 32,
    din309_WIDTH       = 32,
    din310_WIDTH       = 32,
    din311_WIDTH       = 32,
    din312_WIDTH       = 32,
    din313_WIDTH       = 32,
    din314_WIDTH       = 32,
    din315_WIDTH       = 32,
    din316_WIDTH       = 32,
    din317_WIDTH       = 32,
    din318_WIDTH       = 32,
    din319_WIDTH       = 32,
    din320_WIDTH       = 32,
    din321_WIDTH       = 32,
    din322_WIDTH       = 32,
    din323_WIDTH       = 32,
    din324_WIDTH       = 32,
    din325_WIDTH       = 32,
    din326_WIDTH       = 32,
    din327_WIDTH       = 32,
    din328_WIDTH       = 32,
    din329_WIDTH       = 32,
    din330_WIDTH       = 32,
    din331_WIDTH       = 32,
    din332_WIDTH       = 32,
    din333_WIDTH       = 32,
    din334_WIDTH       = 32,
    din335_WIDTH       = 32,
    din336_WIDTH       = 32,
    din337_WIDTH       = 32,
    din338_WIDTH       = 32,
    din339_WIDTH       = 32,
    din340_WIDTH       = 32,
    din341_WIDTH       = 32,
    din342_WIDTH       = 32,
    din343_WIDTH       = 32,
    din344_WIDTH       = 32,
    din345_WIDTH       = 32,
    din346_WIDTH       = 32,
    din347_WIDTH       = 32,
    din348_WIDTH       = 32,
    din349_WIDTH       = 32,
    din350_WIDTH       = 32,
    din351_WIDTH       = 32,
    din352_WIDTH       = 32,
    din353_WIDTH       = 32,
    din354_WIDTH       = 32,
    din355_WIDTH       = 32,
    din356_WIDTH       = 32,
    din357_WIDTH       = 32,
    din358_WIDTH       = 32,
    din359_WIDTH       = 32,
    din360_WIDTH       = 32,
    din361_WIDTH       = 32,
    din362_WIDTH       = 32,
    din363_WIDTH       = 32,
    din364_WIDTH       = 32,
    din365_WIDTH       = 32,
    din366_WIDTH       = 32,
    din367_WIDTH       = 32,
    din368_WIDTH       = 32,
    din369_WIDTH       = 32,
    din370_WIDTH       = 32,
    din371_WIDTH       = 32,
    din372_WIDTH       = 32,
    din373_WIDTH       = 32,
    din374_WIDTH       = 32,
    din375_WIDTH       = 32,
    din376_WIDTH       = 32,
    din377_WIDTH       = 32,
    din378_WIDTH       = 32,
    din379_WIDTH       = 32,
    din380_WIDTH       = 32,
    din381_WIDTH       = 32,
    din382_WIDTH       = 32,
    din383_WIDTH       = 32,
    din384_WIDTH       = 32,
    din385_WIDTH       = 32,
    din386_WIDTH       = 32,
    din387_WIDTH       = 32,
    din388_WIDTH       = 32,
    din389_WIDTH       = 32,
    din390_WIDTH       = 32,
    din391_WIDTH       = 32,
    din392_WIDTH       = 32,
    din393_WIDTH       = 32,
    din394_WIDTH       = 32,
    din395_WIDTH       = 32,
    din396_WIDTH       = 32,
    din397_WIDTH       = 32,
    din398_WIDTH       = 32,
    din399_WIDTH       = 32,
    din400_WIDTH       = 32,
    din401_WIDTH       = 32,
    din402_WIDTH       = 32,
    din403_WIDTH       = 32,
    din404_WIDTH       = 32,
    din405_WIDTH       = 32,
    din406_WIDTH       = 32,
    din407_WIDTH       = 32,
    din408_WIDTH       = 32,
    din409_WIDTH       = 32,
    din410_WIDTH       = 32,
    din411_WIDTH       = 32,
    din412_WIDTH       = 32,
    din413_WIDTH       = 32,
    din414_WIDTH       = 32,
    din415_WIDTH       = 32,
    din416_WIDTH       = 32,
    din417_WIDTH       = 32,
    din418_WIDTH       = 32,
    din419_WIDTH       = 32,
    din420_WIDTH       = 32,
    din421_WIDTH       = 32,
    din422_WIDTH       = 32,
    din423_WIDTH       = 32,
    din424_WIDTH       = 32,
    din425_WIDTH       = 32,
    din426_WIDTH       = 32,
    din427_WIDTH       = 32,
    din428_WIDTH       = 32,
    din429_WIDTH       = 32,
    din430_WIDTH       = 32,
    din431_WIDTH       = 32,
    din432_WIDTH       = 32,
    din433_WIDTH       = 32,
    din434_WIDTH       = 32,
    din435_WIDTH       = 32,
    din436_WIDTH       = 32,
    din437_WIDTH       = 32,
    din438_WIDTH       = 32,
    din439_WIDTH       = 32,
    din440_WIDTH       = 32,
    din441_WIDTH       = 32,
    din442_WIDTH       = 32,
    din443_WIDTH       = 32,
    din444_WIDTH       = 32,
    din445_WIDTH       = 32,
    din446_WIDTH       = 32,
    din447_WIDTH       = 32,
    din448_WIDTH       = 32,
    din449_WIDTH       = 32,
    din450_WIDTH       = 32,
    din451_WIDTH       = 32,
    din452_WIDTH       = 32,
    din453_WIDTH       = 32,
    din454_WIDTH       = 32,
    din455_WIDTH       = 32,
    din456_WIDTH       = 32,
    din457_WIDTH       = 32,
    din458_WIDTH       = 32,
    din459_WIDTH       = 32,
    din460_WIDTH       = 32,
    din461_WIDTH       = 32,
    din462_WIDTH       = 32,
    din463_WIDTH       = 32,
    din464_WIDTH       = 32,
    din465_WIDTH       = 32,
    din466_WIDTH       = 32,
    din467_WIDTH       = 32,
    din468_WIDTH       = 32,
    din469_WIDTH       = 32,
    din470_WIDTH       = 32,
    din471_WIDTH       = 32,
    din472_WIDTH       = 32,
    din473_WIDTH       = 32,
    din474_WIDTH       = 32,
    din475_WIDTH       = 32,
    din476_WIDTH       = 32,
    din477_WIDTH       = 32,
    din478_WIDTH       = 32,
    din479_WIDTH       = 32,
    din480_WIDTH       = 32,
    din481_WIDTH       = 32,
    din482_WIDTH       = 32,
    din483_WIDTH       = 32,
    din484_WIDTH       = 32,
    din485_WIDTH       = 32,
    din486_WIDTH       = 32,
    din487_WIDTH       = 32,
    din488_WIDTH       = 32,
    din489_WIDTH       = 32,
    din490_WIDTH       = 32,
    din491_WIDTH       = 32,
    din492_WIDTH       = 32,
    din493_WIDTH       = 32,
    din494_WIDTH       = 32,
    din495_WIDTH       = 32,
    din496_WIDTH       = 32,
    din497_WIDTH       = 32,
    din498_WIDTH       = 32,
    din499_WIDTH       = 32,
    din500_WIDTH       = 32,
    din501_WIDTH       = 32,
    din502_WIDTH       = 32,
    din503_WIDTH       = 32,
    din504_WIDTH       = 32,
    din505_WIDTH       = 32,
    din506_WIDTH       = 32,
    din507_WIDTH       = 32,
    din508_WIDTH       = 32,
    din509_WIDTH       = 32,
    din510_WIDTH       = 32,
    din511_WIDTH       = 32,
    din512_WIDTH       = 32,
    din513_WIDTH       = 32,
    din514_WIDTH       = 32,
    din515_WIDTH       = 32,
    din516_WIDTH       = 32,
    din517_WIDTH       = 32,
    din518_WIDTH       = 32,
    din519_WIDTH       = 32,
    din520_WIDTH       = 32,
    din521_WIDTH       = 32,
    din522_WIDTH       = 32,
    din523_WIDTH       = 32,
    din524_WIDTH       = 32,
    din525_WIDTH       = 32,
    din526_WIDTH       = 32,
    din527_WIDTH       = 32,
    din528_WIDTH       = 32,
    din529_WIDTH       = 32,
    din530_WIDTH       = 32,
    din531_WIDTH       = 32,
    din532_WIDTH       = 32,
    din533_WIDTH       = 32,
    din534_WIDTH       = 32,
    din535_WIDTH       = 32,
    din536_WIDTH       = 32,
    din537_WIDTH       = 32,
    din538_WIDTH       = 32,
    din539_WIDTH       = 32,
    din540_WIDTH       = 32,
    din541_WIDTH       = 32,
    din542_WIDTH       = 32,
    din543_WIDTH       = 32,
    din544_WIDTH       = 32,
    din545_WIDTH       = 32,
    din546_WIDTH       = 32,
    din547_WIDTH       = 32,
    din548_WIDTH       = 32,
    din549_WIDTH       = 32,
    din550_WIDTH       = 32,
    din551_WIDTH       = 32,
    din552_WIDTH       = 32,
    din553_WIDTH       = 32,
    din554_WIDTH       = 32,
    din555_WIDTH       = 32,
    din556_WIDTH       = 32,
    din557_WIDTH       = 32,
    din558_WIDTH       = 32,
    din559_WIDTH       = 32,
    din560_WIDTH       = 32,
    din561_WIDTH       = 32,
    din562_WIDTH       = 32,
    din563_WIDTH       = 32,
    din564_WIDTH       = 32,
    din565_WIDTH       = 32,
    din566_WIDTH       = 32,
    din567_WIDTH       = 32,
    din568_WIDTH       = 32,
    din569_WIDTH       = 32,
    din570_WIDTH       = 32,
    din571_WIDTH       = 32,
    din572_WIDTH       = 32,
    din573_WIDTH       = 32,
    din574_WIDTH       = 32,
    din575_WIDTH       = 32,
    din576_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [7 : 0]     din0,
    input  [7 : 0]     din1,
    input  [7 : 0]     din2,
    input  [7 : 0]     din3,
    input  [7 : 0]     din4,
    input  [7 : 0]     din5,
    input  [7 : 0]     din6,
    input  [7 : 0]     din7,
    input  [7 : 0]     din8,
    input  [7 : 0]     din9,
    input  [7 : 0]     din10,
    input  [7 : 0]     din11,
    input  [7 : 0]     din12,
    input  [7 : 0]     din13,
    input  [7 : 0]     din14,
    input  [7 : 0]     din15,
    input  [7 : 0]     din16,
    input  [7 : 0]     din17,
    input  [7 : 0]     din18,
    input  [7 : 0]     din19,
    input  [7 : 0]     din20,
    input  [7 : 0]     din21,
    input  [7 : 0]     din22,
    input  [7 : 0]     din23,
    input  [7 : 0]     din24,
    input  [7 : 0]     din25,
    input  [7 : 0]     din26,
    input  [7 : 0]     din27,
    input  [7 : 0]     din28,
    input  [7 : 0]     din29,
    input  [7 : 0]     din30,
    input  [7 : 0]     din31,
    input  [7 : 0]     din32,
    input  [7 : 0]     din33,
    input  [7 : 0]     din34,
    input  [7 : 0]     din35,
    input  [7 : 0]     din36,
    input  [7 : 0]     din37,
    input  [7 : 0]     din38,
    input  [7 : 0]     din39,
    input  [7 : 0]     din40,
    input  [7 : 0]     din41,
    input  [7 : 0]     din42,
    input  [7 : 0]     din43,
    input  [7 : 0]     din44,
    input  [7 : 0]     din45,
    input  [7 : 0]     din46,
    input  [7 : 0]     din47,
    input  [7 : 0]     din48,
    input  [7 : 0]     din49,
    input  [7 : 0]     din50,
    input  [7 : 0]     din51,
    input  [7 : 0]     din52,
    input  [7 : 0]     din53,
    input  [7 : 0]     din54,
    input  [7 : 0]     din55,
    input  [7 : 0]     din56,
    input  [7 : 0]     din57,
    input  [7 : 0]     din58,
    input  [7 : 0]     din59,
    input  [7 : 0]     din60,
    input  [7 : 0]     din61,
    input  [7 : 0]     din62,
    input  [7 : 0]     din63,
    input  [7 : 0]     din64,
    input  [7 : 0]     din65,
    input  [7 : 0]     din66,
    input  [7 : 0]     din67,
    input  [7 : 0]     din68,
    input  [7 : 0]     din69,
    input  [7 : 0]     din70,
    input  [7 : 0]     din71,
    input  [7 : 0]     din72,
    input  [7 : 0]     din73,
    input  [7 : 0]     din74,
    input  [7 : 0]     din75,
    input  [7 : 0]     din76,
    input  [7 : 0]     din77,
    input  [7 : 0]     din78,
    input  [7 : 0]     din79,
    input  [7 : 0]     din80,
    input  [7 : 0]     din81,
    input  [7 : 0]     din82,
    input  [7 : 0]     din83,
    input  [7 : 0]     din84,
    input  [7 : 0]     din85,
    input  [7 : 0]     din86,
    input  [7 : 0]     din87,
    input  [7 : 0]     din88,
    input  [7 : 0]     din89,
    input  [7 : 0]     din90,
    input  [7 : 0]     din91,
    input  [7 : 0]     din92,
    input  [7 : 0]     din93,
    input  [7 : 0]     din94,
    input  [7 : 0]     din95,
    input  [7 : 0]     din96,
    input  [7 : 0]     din97,
    input  [7 : 0]     din98,
    input  [7 : 0]     din99,
    input  [7 : 0]     din100,
    input  [7 : 0]     din101,
    input  [7 : 0]     din102,
    input  [7 : 0]     din103,
    input  [7 : 0]     din104,
    input  [7 : 0]     din105,
    input  [7 : 0]     din106,
    input  [7 : 0]     din107,
    input  [7 : 0]     din108,
    input  [7 : 0]     din109,
    input  [7 : 0]     din110,
    input  [7 : 0]     din111,
    input  [7 : 0]     din112,
    input  [7 : 0]     din113,
    input  [7 : 0]     din114,
    input  [7 : 0]     din115,
    input  [7 : 0]     din116,
    input  [7 : 0]     din117,
    input  [7 : 0]     din118,
    input  [7 : 0]     din119,
    input  [7 : 0]     din120,
    input  [7 : 0]     din121,
    input  [7 : 0]     din122,
    input  [7 : 0]     din123,
    input  [7 : 0]     din124,
    input  [7 : 0]     din125,
    input  [7 : 0]     din126,
    input  [7 : 0]     din127,
    input  [7 : 0]     din128,
    input  [7 : 0]     din129,
    input  [7 : 0]     din130,
    input  [7 : 0]     din131,
    input  [7 : 0]     din132,
    input  [7 : 0]     din133,
    input  [7 : 0]     din134,
    input  [7 : 0]     din135,
    input  [7 : 0]     din136,
    input  [7 : 0]     din137,
    input  [7 : 0]     din138,
    input  [7 : 0]     din139,
    input  [7 : 0]     din140,
    input  [7 : 0]     din141,
    input  [7 : 0]     din142,
    input  [7 : 0]     din143,
    input  [7 : 0]     din144,
    input  [7 : 0]     din145,
    input  [7 : 0]     din146,
    input  [7 : 0]     din147,
    input  [7 : 0]     din148,
    input  [7 : 0]     din149,
    input  [7 : 0]     din150,
    input  [7 : 0]     din151,
    input  [7 : 0]     din152,
    input  [7 : 0]     din153,
    input  [7 : 0]     din154,
    input  [7 : 0]     din155,
    input  [7 : 0]     din156,
    input  [7 : 0]     din157,
    input  [7 : 0]     din158,
    input  [7 : 0]     din159,
    input  [7 : 0]     din160,
    input  [7 : 0]     din161,
    input  [7 : 0]     din162,
    input  [7 : 0]     din163,
    input  [7 : 0]     din164,
    input  [7 : 0]     din165,
    input  [7 : 0]     din166,
    input  [7 : 0]     din167,
    input  [7 : 0]     din168,
    input  [7 : 0]     din169,
    input  [7 : 0]     din170,
    input  [7 : 0]     din171,
    input  [7 : 0]     din172,
    input  [7 : 0]     din173,
    input  [7 : 0]     din174,
    input  [7 : 0]     din175,
    input  [7 : 0]     din176,
    input  [7 : 0]     din177,
    input  [7 : 0]     din178,
    input  [7 : 0]     din179,
    input  [7 : 0]     din180,
    input  [7 : 0]     din181,
    input  [7 : 0]     din182,
    input  [7 : 0]     din183,
    input  [7 : 0]     din184,
    input  [7 : 0]     din185,
    input  [7 : 0]     din186,
    input  [7 : 0]     din187,
    input  [7 : 0]     din188,
    input  [7 : 0]     din189,
    input  [7 : 0]     din190,
    input  [7 : 0]     din191,
    input  [7 : 0]     din192,
    input  [7 : 0]     din193,
    input  [7 : 0]     din194,
    input  [7 : 0]     din195,
    input  [7 : 0]     din196,
    input  [7 : 0]     din197,
    input  [7 : 0]     din198,
    input  [7 : 0]     din199,
    input  [7 : 0]     din200,
    input  [7 : 0]     din201,
    input  [7 : 0]     din202,
    input  [7 : 0]     din203,
    input  [7 : 0]     din204,
    input  [7 : 0]     din205,
    input  [7 : 0]     din206,
    input  [7 : 0]     din207,
    input  [7 : 0]     din208,
    input  [7 : 0]     din209,
    input  [7 : 0]     din210,
    input  [7 : 0]     din211,
    input  [7 : 0]     din212,
    input  [7 : 0]     din213,
    input  [7 : 0]     din214,
    input  [7 : 0]     din215,
    input  [7 : 0]     din216,
    input  [7 : 0]     din217,
    input  [7 : 0]     din218,
    input  [7 : 0]     din219,
    input  [7 : 0]     din220,
    input  [7 : 0]     din221,
    input  [7 : 0]     din222,
    input  [7 : 0]     din223,
    input  [7 : 0]     din224,
    input  [7 : 0]     din225,
    input  [7 : 0]     din226,
    input  [7 : 0]     din227,
    input  [7 : 0]     din228,
    input  [7 : 0]     din229,
    input  [7 : 0]     din230,
    input  [7 : 0]     din231,
    input  [7 : 0]     din232,
    input  [7 : 0]     din233,
    input  [7 : 0]     din234,
    input  [7 : 0]     din235,
    input  [7 : 0]     din236,
    input  [7 : 0]     din237,
    input  [7 : 0]     din238,
    input  [7 : 0]     din239,
    input  [7 : 0]     din240,
    input  [7 : 0]     din241,
    input  [7 : 0]     din242,
    input  [7 : 0]     din243,
    input  [7 : 0]     din244,
    input  [7 : 0]     din245,
    input  [7 : 0]     din246,
    input  [7 : 0]     din247,
    input  [7 : 0]     din248,
    input  [7 : 0]     din249,
    input  [7 : 0]     din250,
    input  [7 : 0]     din251,
    input  [7 : 0]     din252,
    input  [7 : 0]     din253,
    input  [7 : 0]     din254,
    input  [7 : 0]     din255,
    input  [7 : 0]     din256,
    input  [7 : 0]     din257,
    input  [7 : 0]     din258,
    input  [7 : 0]     din259,
    input  [7 : 0]     din260,
    input  [7 : 0]     din261,
    input  [7 : 0]     din262,
    input  [7 : 0]     din263,
    input  [7 : 0]     din264,
    input  [7 : 0]     din265,
    input  [7 : 0]     din266,
    input  [7 : 0]     din267,
    input  [7 : 0]     din268,
    input  [7 : 0]     din269,
    input  [7 : 0]     din270,
    input  [7 : 0]     din271,
    input  [7 : 0]     din272,
    input  [7 : 0]     din273,
    input  [7 : 0]     din274,
    input  [7 : 0]     din275,
    input  [7 : 0]     din276,
    input  [7 : 0]     din277,
    input  [7 : 0]     din278,
    input  [7 : 0]     din279,
    input  [7 : 0]     din280,
    input  [7 : 0]     din281,
    input  [7 : 0]     din282,
    input  [7 : 0]     din283,
    input  [7 : 0]     din284,
    input  [7 : 0]     din285,
    input  [7 : 0]     din286,
    input  [7 : 0]     din287,
    input  [7 : 0]     din288,
    input  [7 : 0]     din289,
    input  [7 : 0]     din290,
    input  [7 : 0]     din291,
    input  [7 : 0]     din292,
    input  [7 : 0]     din293,
    input  [7 : 0]     din294,
    input  [7 : 0]     din295,
    input  [7 : 0]     din296,
    input  [7 : 0]     din297,
    input  [7 : 0]     din298,
    input  [7 : 0]     din299,
    input  [7 : 0]     din300,
    input  [7 : 0]     din301,
    input  [7 : 0]     din302,
    input  [7 : 0]     din303,
    input  [7 : 0]     din304,
    input  [7 : 0]     din305,
    input  [7 : 0]     din306,
    input  [7 : 0]     din307,
    input  [7 : 0]     din308,
    input  [7 : 0]     din309,
    input  [7 : 0]     din310,
    input  [7 : 0]     din311,
    input  [7 : 0]     din312,
    input  [7 : 0]     din313,
    input  [7 : 0]     din314,
    input  [7 : 0]     din315,
    input  [7 : 0]     din316,
    input  [7 : 0]     din317,
    input  [7 : 0]     din318,
    input  [7 : 0]     din319,
    input  [7 : 0]     din320,
    input  [7 : 0]     din321,
    input  [7 : 0]     din322,
    input  [7 : 0]     din323,
    input  [7 : 0]     din324,
    input  [7 : 0]     din325,
    input  [7 : 0]     din326,
    input  [7 : 0]     din327,
    input  [7 : 0]     din328,
    input  [7 : 0]     din329,
    input  [7 : 0]     din330,
    input  [7 : 0]     din331,
    input  [7 : 0]     din332,
    input  [7 : 0]     din333,
    input  [7 : 0]     din334,
    input  [7 : 0]     din335,
    input  [7 : 0]     din336,
    input  [7 : 0]     din337,
    input  [7 : 0]     din338,
    input  [7 : 0]     din339,
    input  [7 : 0]     din340,
    input  [7 : 0]     din341,
    input  [7 : 0]     din342,
    input  [7 : 0]     din343,
    input  [7 : 0]     din344,
    input  [7 : 0]     din345,
    input  [7 : 0]     din346,
    input  [7 : 0]     din347,
    input  [7 : 0]     din348,
    input  [7 : 0]     din349,
    input  [7 : 0]     din350,
    input  [7 : 0]     din351,
    input  [7 : 0]     din352,
    input  [7 : 0]     din353,
    input  [7 : 0]     din354,
    input  [7 : 0]     din355,
    input  [7 : 0]     din356,
    input  [7 : 0]     din357,
    input  [7 : 0]     din358,
    input  [7 : 0]     din359,
    input  [7 : 0]     din360,
    input  [7 : 0]     din361,
    input  [7 : 0]     din362,
    input  [7 : 0]     din363,
    input  [7 : 0]     din364,
    input  [7 : 0]     din365,
    input  [7 : 0]     din366,
    input  [7 : 0]     din367,
    input  [7 : 0]     din368,
    input  [7 : 0]     din369,
    input  [7 : 0]     din370,
    input  [7 : 0]     din371,
    input  [7 : 0]     din372,
    input  [7 : 0]     din373,
    input  [7 : 0]     din374,
    input  [7 : 0]     din375,
    input  [7 : 0]     din376,
    input  [7 : 0]     din377,
    input  [7 : 0]     din378,
    input  [7 : 0]     din379,
    input  [7 : 0]     din380,
    input  [7 : 0]     din381,
    input  [7 : 0]     din382,
    input  [7 : 0]     din383,
    input  [7 : 0]     din384,
    input  [7 : 0]     din385,
    input  [7 : 0]     din386,
    input  [7 : 0]     din387,
    input  [7 : 0]     din388,
    input  [7 : 0]     din389,
    input  [7 : 0]     din390,
    input  [7 : 0]     din391,
    input  [7 : 0]     din392,
    input  [7 : 0]     din393,
    input  [7 : 0]     din394,
    input  [7 : 0]     din395,
    input  [7 : 0]     din396,
    input  [7 : 0]     din397,
    input  [7 : 0]     din398,
    input  [7 : 0]     din399,
    input  [7 : 0]     din400,
    input  [7 : 0]     din401,
    input  [7 : 0]     din402,
    input  [7 : 0]     din403,
    input  [7 : 0]     din404,
    input  [7 : 0]     din405,
    input  [7 : 0]     din406,
    input  [7 : 0]     din407,
    input  [7 : 0]     din408,
    input  [7 : 0]     din409,
    input  [7 : 0]     din410,
    input  [7 : 0]     din411,
    input  [7 : 0]     din412,
    input  [7 : 0]     din413,
    input  [7 : 0]     din414,
    input  [7 : 0]     din415,
    input  [7 : 0]     din416,
    input  [7 : 0]     din417,
    input  [7 : 0]     din418,
    input  [7 : 0]     din419,
    input  [7 : 0]     din420,
    input  [7 : 0]     din421,
    input  [7 : 0]     din422,
    input  [7 : 0]     din423,
    input  [7 : 0]     din424,
    input  [7 : 0]     din425,
    input  [7 : 0]     din426,
    input  [7 : 0]     din427,
    input  [7 : 0]     din428,
    input  [7 : 0]     din429,
    input  [7 : 0]     din430,
    input  [7 : 0]     din431,
    input  [7 : 0]     din432,
    input  [7 : 0]     din433,
    input  [7 : 0]     din434,
    input  [7 : 0]     din435,
    input  [7 : 0]     din436,
    input  [7 : 0]     din437,
    input  [7 : 0]     din438,
    input  [7 : 0]     din439,
    input  [7 : 0]     din440,
    input  [7 : 0]     din441,
    input  [7 : 0]     din442,
    input  [7 : 0]     din443,
    input  [7 : 0]     din444,
    input  [7 : 0]     din445,
    input  [7 : 0]     din446,
    input  [7 : 0]     din447,
    input  [7 : 0]     din448,
    input  [7 : 0]     din449,
    input  [7 : 0]     din450,
    input  [7 : 0]     din451,
    input  [7 : 0]     din452,
    input  [7 : 0]     din453,
    input  [7 : 0]     din454,
    input  [7 : 0]     din455,
    input  [7 : 0]     din456,
    input  [7 : 0]     din457,
    input  [7 : 0]     din458,
    input  [7 : 0]     din459,
    input  [7 : 0]     din460,
    input  [7 : 0]     din461,
    input  [7 : 0]     din462,
    input  [7 : 0]     din463,
    input  [7 : 0]     din464,
    input  [7 : 0]     din465,
    input  [7 : 0]     din466,
    input  [7 : 0]     din467,
    input  [7 : 0]     din468,
    input  [7 : 0]     din469,
    input  [7 : 0]     din470,
    input  [7 : 0]     din471,
    input  [7 : 0]     din472,
    input  [7 : 0]     din473,
    input  [7 : 0]     din474,
    input  [7 : 0]     din475,
    input  [7 : 0]     din476,
    input  [7 : 0]     din477,
    input  [7 : 0]     din478,
    input  [7 : 0]     din479,
    input  [7 : 0]     din480,
    input  [7 : 0]     din481,
    input  [7 : 0]     din482,
    input  [7 : 0]     din483,
    input  [7 : 0]     din484,
    input  [7 : 0]     din485,
    input  [7 : 0]     din486,
    input  [7 : 0]     din487,
    input  [7 : 0]     din488,
    input  [7 : 0]     din489,
    input  [7 : 0]     din490,
    input  [7 : 0]     din491,
    input  [7 : 0]     din492,
    input  [7 : 0]     din493,
    input  [7 : 0]     din494,
    input  [7 : 0]     din495,
    input  [7 : 0]     din496,
    input  [7 : 0]     din497,
    input  [7 : 0]     din498,
    input  [7 : 0]     din499,
    input  [7 : 0]     din500,
    input  [7 : 0]     din501,
    input  [7 : 0]     din502,
    input  [7 : 0]     din503,
    input  [7 : 0]     din504,
    input  [7 : 0]     din505,
    input  [7 : 0]     din506,
    input  [7 : 0]     din507,
    input  [7 : 0]     din508,
    input  [7 : 0]     din509,
    input  [7 : 0]     din510,
    input  [7 : 0]     din511,
    input  [7 : 0]     din512,
    input  [7 : 0]     din513,
    input  [7 : 0]     din514,
    input  [7 : 0]     din515,
    input  [7 : 0]     din516,
    input  [7 : 0]     din517,
    input  [7 : 0]     din518,
    input  [7 : 0]     din519,
    input  [7 : 0]     din520,
    input  [7 : 0]     din521,
    input  [7 : 0]     din522,
    input  [7 : 0]     din523,
    input  [7 : 0]     din524,
    input  [7 : 0]     din525,
    input  [7 : 0]     din526,
    input  [7 : 0]     din527,
    input  [7 : 0]     din528,
    input  [7 : 0]     din529,
    input  [7 : 0]     din530,
    input  [7 : 0]     din531,
    input  [7 : 0]     din532,
    input  [7 : 0]     din533,
    input  [7 : 0]     din534,
    input  [7 : 0]     din535,
    input  [7 : 0]     din536,
    input  [7 : 0]     din537,
    input  [7 : 0]     din538,
    input  [7 : 0]     din539,
    input  [7 : 0]     din540,
    input  [7 : 0]     din541,
    input  [7 : 0]     din542,
    input  [7 : 0]     din543,
    input  [7 : 0]     din544,
    input  [7 : 0]     din545,
    input  [7 : 0]     din546,
    input  [7 : 0]     din547,
    input  [7 : 0]     din548,
    input  [7 : 0]     din549,
    input  [7 : 0]     din550,
    input  [7 : 0]     din551,
    input  [7 : 0]     din552,
    input  [7 : 0]     din553,
    input  [7 : 0]     din554,
    input  [7 : 0]     din555,
    input  [7 : 0]     din556,
    input  [7 : 0]     din557,
    input  [7 : 0]     din558,
    input  [7 : 0]     din559,
    input  [7 : 0]     din560,
    input  [7 : 0]     din561,
    input  [7 : 0]     din562,
    input  [7 : 0]     din563,
    input  [7 : 0]     din564,
    input  [7 : 0]     din565,
    input  [7 : 0]     din566,
    input  [7 : 0]     din567,
    input  [7 : 0]     din568,
    input  [7 : 0]     din569,
    input  [7 : 0]     din570,
    input  [7 : 0]     din571,
    input  [7 : 0]     din572,
    input  [7 : 0]     din573,
    input  [7 : 0]     din574,
    input  [7 : 0]     din575,
    input  [9 : 0]    din576,
    output [7 : 0]   dout);

// puts internal signals
wire [9 : 0]     sel;
// level 1 signals
wire [7 : 0]         mux_1_0;
wire [7 : 0]         mux_1_1;
wire [7 : 0]         mux_1_2;
wire [7 : 0]         mux_1_3;
wire [7 : 0]         mux_1_4;
wire [7 : 0]         mux_1_5;
wire [7 : 0]         mux_1_6;
wire [7 : 0]         mux_1_7;
wire [7 : 0]         mux_1_8;
wire [7 : 0]         mux_1_9;
wire [7 : 0]         mux_1_10;
wire [7 : 0]         mux_1_11;
wire [7 : 0]         mux_1_12;
wire [7 : 0]         mux_1_13;
wire [7 : 0]         mux_1_14;
wire [7 : 0]         mux_1_15;
wire [7 : 0]         mux_1_16;
wire [7 : 0]         mux_1_17;
wire [7 : 0]         mux_1_18;
wire [7 : 0]         mux_1_19;
wire [7 : 0]         mux_1_20;
wire [7 : 0]         mux_1_21;
wire [7 : 0]         mux_1_22;
wire [7 : 0]         mux_1_23;
wire [7 : 0]         mux_1_24;
wire [7 : 0]         mux_1_25;
wire [7 : 0]         mux_1_26;
wire [7 : 0]         mux_1_27;
wire [7 : 0]         mux_1_28;
wire [7 : 0]         mux_1_29;
wire [7 : 0]         mux_1_30;
wire [7 : 0]         mux_1_31;
wire [7 : 0]         mux_1_32;
wire [7 : 0]         mux_1_33;
wire [7 : 0]         mux_1_34;
wire [7 : 0]         mux_1_35;
wire [7 : 0]         mux_1_36;
wire [7 : 0]         mux_1_37;
wire [7 : 0]         mux_1_38;
wire [7 : 0]         mux_1_39;
wire [7 : 0]         mux_1_40;
wire [7 : 0]         mux_1_41;
wire [7 : 0]         mux_1_42;
wire [7 : 0]         mux_1_43;
wire [7 : 0]         mux_1_44;
wire [7 : 0]         mux_1_45;
wire [7 : 0]         mux_1_46;
wire [7 : 0]         mux_1_47;
wire [7 : 0]         mux_1_48;
wire [7 : 0]         mux_1_49;
wire [7 : 0]         mux_1_50;
wire [7 : 0]         mux_1_51;
wire [7 : 0]         mux_1_52;
wire [7 : 0]         mux_1_53;
wire [7 : 0]         mux_1_54;
wire [7 : 0]         mux_1_55;
wire [7 : 0]         mux_1_56;
wire [7 : 0]         mux_1_57;
wire [7 : 0]         mux_1_58;
wire [7 : 0]         mux_1_59;
wire [7 : 0]         mux_1_60;
wire [7 : 0]         mux_1_61;
wire [7 : 0]         mux_1_62;
wire [7 : 0]         mux_1_63;
wire [7 : 0]         mux_1_64;
wire [7 : 0]         mux_1_65;
wire [7 : 0]         mux_1_66;
wire [7 : 0]         mux_1_67;
wire [7 : 0]         mux_1_68;
wire [7 : 0]         mux_1_69;
wire [7 : 0]         mux_1_70;
wire [7 : 0]         mux_1_71;
wire [7 : 0]         mux_1_72;
wire [7 : 0]         mux_1_73;
wire [7 : 0]         mux_1_74;
wire [7 : 0]         mux_1_75;
wire [7 : 0]         mux_1_76;
wire [7 : 0]         mux_1_77;
wire [7 : 0]         mux_1_78;
wire [7 : 0]         mux_1_79;
wire [7 : 0]         mux_1_80;
wire [7 : 0]         mux_1_81;
wire [7 : 0]         mux_1_82;
wire [7 : 0]         mux_1_83;
wire [7 : 0]         mux_1_84;
wire [7 : 0]         mux_1_85;
wire [7 : 0]         mux_1_86;
wire [7 : 0]         mux_1_87;
wire [7 : 0]         mux_1_88;
wire [7 : 0]         mux_1_89;
wire [7 : 0]         mux_1_90;
wire [7 : 0]         mux_1_91;
wire [7 : 0]         mux_1_92;
wire [7 : 0]         mux_1_93;
wire [7 : 0]         mux_1_94;
wire [7 : 0]         mux_1_95;
wire [7 : 0]         mux_1_96;
wire [7 : 0]         mux_1_97;
wire [7 : 0]         mux_1_98;
wire [7 : 0]         mux_1_99;
wire [7 : 0]         mux_1_100;
wire [7 : 0]         mux_1_101;
wire [7 : 0]         mux_1_102;
wire [7 : 0]         mux_1_103;
wire [7 : 0]         mux_1_104;
wire [7 : 0]         mux_1_105;
wire [7 : 0]         mux_1_106;
wire [7 : 0]         mux_1_107;
wire [7 : 0]         mux_1_108;
wire [7 : 0]         mux_1_109;
wire [7 : 0]         mux_1_110;
wire [7 : 0]         mux_1_111;
wire [7 : 0]         mux_1_112;
wire [7 : 0]         mux_1_113;
wire [7 : 0]         mux_1_114;
wire [7 : 0]         mux_1_115;
wire [7 : 0]         mux_1_116;
wire [7 : 0]         mux_1_117;
wire [7 : 0]         mux_1_118;
wire [7 : 0]         mux_1_119;
wire [7 : 0]         mux_1_120;
wire [7 : 0]         mux_1_121;
wire [7 : 0]         mux_1_122;
wire [7 : 0]         mux_1_123;
wire [7 : 0]         mux_1_124;
wire [7 : 0]         mux_1_125;
wire [7 : 0]         mux_1_126;
wire [7 : 0]         mux_1_127;
wire [7 : 0]         mux_1_128;
wire [7 : 0]         mux_1_129;
wire [7 : 0]         mux_1_130;
wire [7 : 0]         mux_1_131;
wire [7 : 0]         mux_1_132;
wire [7 : 0]         mux_1_133;
wire [7 : 0]         mux_1_134;
wire [7 : 0]         mux_1_135;
wire [7 : 0]         mux_1_136;
wire [7 : 0]         mux_1_137;
wire [7 : 0]         mux_1_138;
wire [7 : 0]         mux_1_139;
wire [7 : 0]         mux_1_140;
wire [7 : 0]         mux_1_141;
wire [7 : 0]         mux_1_142;
wire [7 : 0]         mux_1_143;
wire [7 : 0]         mux_1_144;
wire [7 : 0]         mux_1_145;
wire [7 : 0]         mux_1_146;
wire [7 : 0]         mux_1_147;
wire [7 : 0]         mux_1_148;
wire [7 : 0]         mux_1_149;
wire [7 : 0]         mux_1_150;
wire [7 : 0]         mux_1_151;
wire [7 : 0]         mux_1_152;
wire [7 : 0]         mux_1_153;
wire [7 : 0]         mux_1_154;
wire [7 : 0]         mux_1_155;
wire [7 : 0]         mux_1_156;
wire [7 : 0]         mux_1_157;
wire [7 : 0]         mux_1_158;
wire [7 : 0]         mux_1_159;
wire [7 : 0]         mux_1_160;
wire [7 : 0]         mux_1_161;
wire [7 : 0]         mux_1_162;
wire [7 : 0]         mux_1_163;
wire [7 : 0]         mux_1_164;
wire [7 : 0]         mux_1_165;
wire [7 : 0]         mux_1_166;
wire [7 : 0]         mux_1_167;
wire [7 : 0]         mux_1_168;
wire [7 : 0]         mux_1_169;
wire [7 : 0]         mux_1_170;
wire [7 : 0]         mux_1_171;
wire [7 : 0]         mux_1_172;
wire [7 : 0]         mux_1_173;
wire [7 : 0]         mux_1_174;
wire [7 : 0]         mux_1_175;
wire [7 : 0]         mux_1_176;
wire [7 : 0]         mux_1_177;
wire [7 : 0]         mux_1_178;
wire [7 : 0]         mux_1_179;
wire [7 : 0]         mux_1_180;
wire [7 : 0]         mux_1_181;
wire [7 : 0]         mux_1_182;
wire [7 : 0]         mux_1_183;
wire [7 : 0]         mux_1_184;
wire [7 : 0]         mux_1_185;
wire [7 : 0]         mux_1_186;
wire [7 : 0]         mux_1_187;
wire [7 : 0]         mux_1_188;
wire [7 : 0]         mux_1_189;
wire [7 : 0]         mux_1_190;
wire [7 : 0]         mux_1_191;
wire [7 : 0]         mux_1_192;
wire [7 : 0]         mux_1_193;
wire [7 : 0]         mux_1_194;
wire [7 : 0]         mux_1_195;
wire [7 : 0]         mux_1_196;
wire [7 : 0]         mux_1_197;
wire [7 : 0]         mux_1_198;
wire [7 : 0]         mux_1_199;
wire [7 : 0]         mux_1_200;
wire [7 : 0]         mux_1_201;
wire [7 : 0]         mux_1_202;
wire [7 : 0]         mux_1_203;
wire [7 : 0]         mux_1_204;
wire [7 : 0]         mux_1_205;
wire [7 : 0]         mux_1_206;
wire [7 : 0]         mux_1_207;
wire [7 : 0]         mux_1_208;
wire [7 : 0]         mux_1_209;
wire [7 : 0]         mux_1_210;
wire [7 : 0]         mux_1_211;
wire [7 : 0]         mux_1_212;
wire [7 : 0]         mux_1_213;
wire [7 : 0]         mux_1_214;
wire [7 : 0]         mux_1_215;
wire [7 : 0]         mux_1_216;
wire [7 : 0]         mux_1_217;
wire [7 : 0]         mux_1_218;
wire [7 : 0]         mux_1_219;
wire [7 : 0]         mux_1_220;
wire [7 : 0]         mux_1_221;
wire [7 : 0]         mux_1_222;
wire [7 : 0]         mux_1_223;
wire [7 : 0]         mux_1_224;
wire [7 : 0]         mux_1_225;
wire [7 : 0]         mux_1_226;
wire [7 : 0]         mux_1_227;
wire [7 : 0]         mux_1_228;
wire [7 : 0]         mux_1_229;
wire [7 : 0]         mux_1_230;
wire [7 : 0]         mux_1_231;
wire [7 : 0]         mux_1_232;
wire [7 : 0]         mux_1_233;
wire [7 : 0]         mux_1_234;
wire [7 : 0]         mux_1_235;
wire [7 : 0]         mux_1_236;
wire [7 : 0]         mux_1_237;
wire [7 : 0]         mux_1_238;
wire [7 : 0]         mux_1_239;
wire [7 : 0]         mux_1_240;
wire [7 : 0]         mux_1_241;
wire [7 : 0]         mux_1_242;
wire [7 : 0]         mux_1_243;
wire [7 : 0]         mux_1_244;
wire [7 : 0]         mux_1_245;
wire [7 : 0]         mux_1_246;
wire [7 : 0]         mux_1_247;
wire [7 : 0]         mux_1_248;
wire [7 : 0]         mux_1_249;
wire [7 : 0]         mux_1_250;
wire [7 : 0]         mux_1_251;
wire [7 : 0]         mux_1_252;
wire [7 : 0]         mux_1_253;
wire [7 : 0]         mux_1_254;
wire [7 : 0]         mux_1_255;
wire [7 : 0]         mux_1_256;
wire [7 : 0]         mux_1_257;
wire [7 : 0]         mux_1_258;
wire [7 : 0]         mux_1_259;
wire [7 : 0]         mux_1_260;
wire [7 : 0]         mux_1_261;
wire [7 : 0]         mux_1_262;
wire [7 : 0]         mux_1_263;
wire [7 : 0]         mux_1_264;
wire [7 : 0]         mux_1_265;
wire [7 : 0]         mux_1_266;
wire [7 : 0]         mux_1_267;
wire [7 : 0]         mux_1_268;
wire [7 : 0]         mux_1_269;
wire [7 : 0]         mux_1_270;
wire [7 : 0]         mux_1_271;
wire [7 : 0]         mux_1_272;
wire [7 : 0]         mux_1_273;
wire [7 : 0]         mux_1_274;
wire [7 : 0]         mux_1_275;
wire [7 : 0]         mux_1_276;
wire [7 : 0]         mux_1_277;
wire [7 : 0]         mux_1_278;
wire [7 : 0]         mux_1_279;
wire [7 : 0]         mux_1_280;
wire [7 : 0]         mux_1_281;
wire [7 : 0]         mux_1_282;
wire [7 : 0]         mux_1_283;
wire [7 : 0]         mux_1_284;
wire [7 : 0]         mux_1_285;
wire [7 : 0]         mux_1_286;
wire [7 : 0]         mux_1_287;
// level 2 signals
wire [7 : 0]         mux_2_0;
wire [7 : 0]         mux_2_1;
wire [7 : 0]         mux_2_2;
wire [7 : 0]         mux_2_3;
wire [7 : 0]         mux_2_4;
wire [7 : 0]         mux_2_5;
wire [7 : 0]         mux_2_6;
wire [7 : 0]         mux_2_7;
wire [7 : 0]         mux_2_8;
wire [7 : 0]         mux_2_9;
wire [7 : 0]         mux_2_10;
wire [7 : 0]         mux_2_11;
wire [7 : 0]         mux_2_12;
wire [7 : 0]         mux_2_13;
wire [7 : 0]         mux_2_14;
wire [7 : 0]         mux_2_15;
wire [7 : 0]         mux_2_16;
wire [7 : 0]         mux_2_17;
wire [7 : 0]         mux_2_18;
wire [7 : 0]         mux_2_19;
wire [7 : 0]         mux_2_20;
wire [7 : 0]         mux_2_21;
wire [7 : 0]         mux_2_22;
wire [7 : 0]         mux_2_23;
wire [7 : 0]         mux_2_24;
wire [7 : 0]         mux_2_25;
wire [7 : 0]         mux_2_26;
wire [7 : 0]         mux_2_27;
wire [7 : 0]         mux_2_28;
wire [7 : 0]         mux_2_29;
wire [7 : 0]         mux_2_30;
wire [7 : 0]         mux_2_31;
wire [7 : 0]         mux_2_32;
wire [7 : 0]         mux_2_33;
wire [7 : 0]         mux_2_34;
wire [7 : 0]         mux_2_35;
wire [7 : 0]         mux_2_36;
wire [7 : 0]         mux_2_37;
wire [7 : 0]         mux_2_38;
wire [7 : 0]         mux_2_39;
wire [7 : 0]         mux_2_40;
wire [7 : 0]         mux_2_41;
wire [7 : 0]         mux_2_42;
wire [7 : 0]         mux_2_43;
wire [7 : 0]         mux_2_44;
wire [7 : 0]         mux_2_45;
wire [7 : 0]         mux_2_46;
wire [7 : 0]         mux_2_47;
wire [7 : 0]         mux_2_48;
wire [7 : 0]         mux_2_49;
wire [7 : 0]         mux_2_50;
wire [7 : 0]         mux_2_51;
wire [7 : 0]         mux_2_52;
wire [7 : 0]         mux_2_53;
wire [7 : 0]         mux_2_54;
wire [7 : 0]         mux_2_55;
wire [7 : 0]         mux_2_56;
wire [7 : 0]         mux_2_57;
wire [7 : 0]         mux_2_58;
wire [7 : 0]         mux_2_59;
wire [7 : 0]         mux_2_60;
wire [7 : 0]         mux_2_61;
wire [7 : 0]         mux_2_62;
wire [7 : 0]         mux_2_63;
wire [7 : 0]         mux_2_64;
wire [7 : 0]         mux_2_65;
wire [7 : 0]         mux_2_66;
wire [7 : 0]         mux_2_67;
wire [7 : 0]         mux_2_68;
wire [7 : 0]         mux_2_69;
wire [7 : 0]         mux_2_70;
wire [7 : 0]         mux_2_71;
wire [7 : 0]         mux_2_72;
wire [7 : 0]         mux_2_73;
wire [7 : 0]         mux_2_74;
wire [7 : 0]         mux_2_75;
wire [7 : 0]         mux_2_76;
wire [7 : 0]         mux_2_77;
wire [7 : 0]         mux_2_78;
wire [7 : 0]         mux_2_79;
wire [7 : 0]         mux_2_80;
wire [7 : 0]         mux_2_81;
wire [7 : 0]         mux_2_82;
wire [7 : 0]         mux_2_83;
wire [7 : 0]         mux_2_84;
wire [7 : 0]         mux_2_85;
wire [7 : 0]         mux_2_86;
wire [7 : 0]         mux_2_87;
wire [7 : 0]         mux_2_88;
wire [7 : 0]         mux_2_89;
wire [7 : 0]         mux_2_90;
wire [7 : 0]         mux_2_91;
wire [7 : 0]         mux_2_92;
wire [7 : 0]         mux_2_93;
wire [7 : 0]         mux_2_94;
wire [7 : 0]         mux_2_95;
wire [7 : 0]         mux_2_96;
wire [7 : 0]         mux_2_97;
wire [7 : 0]         mux_2_98;
wire [7 : 0]         mux_2_99;
wire [7 : 0]         mux_2_100;
wire [7 : 0]         mux_2_101;
wire [7 : 0]         mux_2_102;
wire [7 : 0]         mux_2_103;
wire [7 : 0]         mux_2_104;
wire [7 : 0]         mux_2_105;
wire [7 : 0]         mux_2_106;
wire [7 : 0]         mux_2_107;
wire [7 : 0]         mux_2_108;
wire [7 : 0]         mux_2_109;
wire [7 : 0]         mux_2_110;
wire [7 : 0]         mux_2_111;
wire [7 : 0]         mux_2_112;
wire [7 : 0]         mux_2_113;
wire [7 : 0]         mux_2_114;
wire [7 : 0]         mux_2_115;
wire [7 : 0]         mux_2_116;
wire [7 : 0]         mux_2_117;
wire [7 : 0]         mux_2_118;
wire [7 : 0]         mux_2_119;
wire [7 : 0]         mux_2_120;
wire [7 : 0]         mux_2_121;
wire [7 : 0]         mux_2_122;
wire [7 : 0]         mux_2_123;
wire [7 : 0]         mux_2_124;
wire [7 : 0]         mux_2_125;
wire [7 : 0]         mux_2_126;
wire [7 : 0]         mux_2_127;
wire [7 : 0]         mux_2_128;
wire [7 : 0]         mux_2_129;
wire [7 : 0]         mux_2_130;
wire [7 : 0]         mux_2_131;
wire [7 : 0]         mux_2_132;
wire [7 : 0]         mux_2_133;
wire [7 : 0]         mux_2_134;
wire [7 : 0]         mux_2_135;
wire [7 : 0]         mux_2_136;
wire [7 : 0]         mux_2_137;
wire [7 : 0]         mux_2_138;
wire [7 : 0]         mux_2_139;
wire [7 : 0]         mux_2_140;
wire [7 : 0]         mux_2_141;
wire [7 : 0]         mux_2_142;
wire [7 : 0]         mux_2_143;
// level 3 signals
wire [7 : 0]         mux_3_0;
wire [7 : 0]         mux_3_1;
wire [7 : 0]         mux_3_2;
wire [7 : 0]         mux_3_3;
wire [7 : 0]         mux_3_4;
wire [7 : 0]         mux_3_5;
wire [7 : 0]         mux_3_6;
wire [7 : 0]         mux_3_7;
wire [7 : 0]         mux_3_8;
wire [7 : 0]         mux_3_9;
wire [7 : 0]         mux_3_10;
wire [7 : 0]         mux_3_11;
wire [7 : 0]         mux_3_12;
wire [7 : 0]         mux_3_13;
wire [7 : 0]         mux_3_14;
wire [7 : 0]         mux_3_15;
wire [7 : 0]         mux_3_16;
wire [7 : 0]         mux_3_17;
wire [7 : 0]         mux_3_18;
wire [7 : 0]         mux_3_19;
wire [7 : 0]         mux_3_20;
wire [7 : 0]         mux_3_21;
wire [7 : 0]         mux_3_22;
wire [7 : 0]         mux_3_23;
wire [7 : 0]         mux_3_24;
wire [7 : 0]         mux_3_25;
wire [7 : 0]         mux_3_26;
wire [7 : 0]         mux_3_27;
wire [7 : 0]         mux_3_28;
wire [7 : 0]         mux_3_29;
wire [7 : 0]         mux_3_30;
wire [7 : 0]         mux_3_31;
wire [7 : 0]         mux_3_32;
wire [7 : 0]         mux_3_33;
wire [7 : 0]         mux_3_34;
wire [7 : 0]         mux_3_35;
wire [7 : 0]         mux_3_36;
wire [7 : 0]         mux_3_37;
wire [7 : 0]         mux_3_38;
wire [7 : 0]         mux_3_39;
wire [7 : 0]         mux_3_40;
wire [7 : 0]         mux_3_41;
wire [7 : 0]         mux_3_42;
wire [7 : 0]         mux_3_43;
wire [7 : 0]         mux_3_44;
wire [7 : 0]         mux_3_45;
wire [7 : 0]         mux_3_46;
wire [7 : 0]         mux_3_47;
wire [7 : 0]         mux_3_48;
wire [7 : 0]         mux_3_49;
wire [7 : 0]         mux_3_50;
wire [7 : 0]         mux_3_51;
wire [7 : 0]         mux_3_52;
wire [7 : 0]         mux_3_53;
wire [7 : 0]         mux_3_54;
wire [7 : 0]         mux_3_55;
wire [7 : 0]         mux_3_56;
wire [7 : 0]         mux_3_57;
wire [7 : 0]         mux_3_58;
wire [7 : 0]         mux_3_59;
wire [7 : 0]         mux_3_60;
wire [7 : 0]         mux_3_61;
wire [7 : 0]         mux_3_62;
wire [7 : 0]         mux_3_63;
wire [7 : 0]         mux_3_64;
wire [7 : 0]         mux_3_65;
wire [7 : 0]         mux_3_66;
wire [7 : 0]         mux_3_67;
wire [7 : 0]         mux_3_68;
wire [7 : 0]         mux_3_69;
wire [7 : 0]         mux_3_70;
wire [7 : 0]         mux_3_71;
// level 4 signals
wire [7 : 0]         mux_4_0;
wire [7 : 0]         mux_4_1;
wire [7 : 0]         mux_4_2;
wire [7 : 0]         mux_4_3;
wire [7 : 0]         mux_4_4;
wire [7 : 0]         mux_4_5;
wire [7 : 0]         mux_4_6;
wire [7 : 0]         mux_4_7;
wire [7 : 0]         mux_4_8;
wire [7 : 0]         mux_4_9;
wire [7 : 0]         mux_4_10;
wire [7 : 0]         mux_4_11;
wire [7 : 0]         mux_4_12;
wire [7 : 0]         mux_4_13;
wire [7 : 0]         mux_4_14;
wire [7 : 0]         mux_4_15;
wire [7 : 0]         mux_4_16;
wire [7 : 0]         mux_4_17;
wire [7 : 0]         mux_4_18;
wire [7 : 0]         mux_4_19;
wire [7 : 0]         mux_4_20;
wire [7 : 0]         mux_4_21;
wire [7 : 0]         mux_4_22;
wire [7 : 0]         mux_4_23;
wire [7 : 0]         mux_4_24;
wire [7 : 0]         mux_4_25;
wire [7 : 0]         mux_4_26;
wire [7 : 0]         mux_4_27;
wire [7 : 0]         mux_4_28;
wire [7 : 0]         mux_4_29;
wire [7 : 0]         mux_4_30;
wire [7 : 0]         mux_4_31;
wire [7 : 0]         mux_4_32;
wire [7 : 0]         mux_4_33;
wire [7 : 0]         mux_4_34;
wire [7 : 0]         mux_4_35;
// level 5 signals
wire [7 : 0]         mux_5_0;
wire [7 : 0]         mux_5_1;
wire [7 : 0]         mux_5_2;
wire [7 : 0]         mux_5_3;
wire [7 : 0]         mux_5_4;
wire [7 : 0]         mux_5_5;
wire [7 : 0]         mux_5_6;
wire [7 : 0]         mux_5_7;
wire [7 : 0]         mux_5_8;
wire [7 : 0]         mux_5_9;
wire [7 : 0]         mux_5_10;
wire [7 : 0]         mux_5_11;
wire [7 : 0]         mux_5_12;
wire [7 : 0]         mux_5_13;
wire [7 : 0]         mux_5_14;
wire [7 : 0]         mux_5_15;
wire [7 : 0]         mux_5_16;
wire [7 : 0]         mux_5_17;
// level 6 signals
wire [7 : 0]         mux_6_0;
wire [7 : 0]         mux_6_1;
wire [7 : 0]         mux_6_2;
wire [7 : 0]         mux_6_3;
wire [7 : 0]         mux_6_4;
wire [7 : 0]         mux_6_5;
wire [7 : 0]         mux_6_6;
wire [7 : 0]         mux_6_7;
wire [7 : 0]         mux_6_8;
// level 7 signals
wire [7 : 0]         mux_7_0;
wire [7 : 0]         mux_7_1;
wire [7 : 0]         mux_7_2;
wire [7 : 0]         mux_7_3;
wire [7 : 0]         mux_7_4;
// level 8 signals
wire [7 : 0]         mux_8_0;
wire [7 : 0]         mux_8_1;
wire [7 : 0]         mux_8_2;
// level 9 signals
wire [7 : 0]         mux_9_0;
wire [7 : 0]         mux_9_1;
// level 10 signals
wire [7 : 0]         mux_10_0;

assign sel = din576;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;
assign mux_1_2 = (sel[0] == 0)? din4 : din5;
assign mux_1_3 = (sel[0] == 0)? din6 : din7;
assign mux_1_4 = (sel[0] == 0)? din8 : din9;
assign mux_1_5 = (sel[0] == 0)? din10 : din11;
assign mux_1_6 = (sel[0] == 0)? din12 : din13;
assign mux_1_7 = (sel[0] == 0)? din14 : din15;
assign mux_1_8 = (sel[0] == 0)? din16 : din17;
assign mux_1_9 = (sel[0] == 0)? din18 : din19;
assign mux_1_10 = (sel[0] == 0)? din20 : din21;
assign mux_1_11 = (sel[0] == 0)? din22 : din23;
assign mux_1_12 = (sel[0] == 0)? din24 : din25;
assign mux_1_13 = (sel[0] == 0)? din26 : din27;
assign mux_1_14 = (sel[0] == 0)? din28 : din29;
assign mux_1_15 = (sel[0] == 0)? din30 : din31;
assign mux_1_16 = (sel[0] == 0)? din32 : din33;
assign mux_1_17 = (sel[0] == 0)? din34 : din35;
assign mux_1_18 = (sel[0] == 0)? din36 : din37;
assign mux_1_19 = (sel[0] == 0)? din38 : din39;
assign mux_1_20 = (sel[0] == 0)? din40 : din41;
assign mux_1_21 = (sel[0] == 0)? din42 : din43;
assign mux_1_22 = (sel[0] == 0)? din44 : din45;
assign mux_1_23 = (sel[0] == 0)? din46 : din47;
assign mux_1_24 = (sel[0] == 0)? din48 : din49;
assign mux_1_25 = (sel[0] == 0)? din50 : din51;
assign mux_1_26 = (sel[0] == 0)? din52 : din53;
assign mux_1_27 = (sel[0] == 0)? din54 : din55;
assign mux_1_28 = (sel[0] == 0)? din56 : din57;
assign mux_1_29 = (sel[0] == 0)? din58 : din59;
assign mux_1_30 = (sel[0] == 0)? din60 : din61;
assign mux_1_31 = (sel[0] == 0)? din62 : din63;
assign mux_1_32 = (sel[0] == 0)? din64 : din65;
assign mux_1_33 = (sel[0] == 0)? din66 : din67;
assign mux_1_34 = (sel[0] == 0)? din68 : din69;
assign mux_1_35 = (sel[0] == 0)? din70 : din71;
assign mux_1_36 = (sel[0] == 0)? din72 : din73;
assign mux_1_37 = (sel[0] == 0)? din74 : din75;
assign mux_1_38 = (sel[0] == 0)? din76 : din77;
assign mux_1_39 = (sel[0] == 0)? din78 : din79;
assign mux_1_40 = (sel[0] == 0)? din80 : din81;
assign mux_1_41 = (sel[0] == 0)? din82 : din83;
assign mux_1_42 = (sel[0] == 0)? din84 : din85;
assign mux_1_43 = (sel[0] == 0)? din86 : din87;
assign mux_1_44 = (sel[0] == 0)? din88 : din89;
assign mux_1_45 = (sel[0] == 0)? din90 : din91;
assign mux_1_46 = (sel[0] == 0)? din92 : din93;
assign mux_1_47 = (sel[0] == 0)? din94 : din95;
assign mux_1_48 = (sel[0] == 0)? din96 : din97;
assign mux_1_49 = (sel[0] == 0)? din98 : din99;
assign mux_1_50 = (sel[0] == 0)? din100 : din101;
assign mux_1_51 = (sel[0] == 0)? din102 : din103;
assign mux_1_52 = (sel[0] == 0)? din104 : din105;
assign mux_1_53 = (sel[0] == 0)? din106 : din107;
assign mux_1_54 = (sel[0] == 0)? din108 : din109;
assign mux_1_55 = (sel[0] == 0)? din110 : din111;
assign mux_1_56 = (sel[0] == 0)? din112 : din113;
assign mux_1_57 = (sel[0] == 0)? din114 : din115;
assign mux_1_58 = (sel[0] == 0)? din116 : din117;
assign mux_1_59 = (sel[0] == 0)? din118 : din119;
assign mux_1_60 = (sel[0] == 0)? din120 : din121;
assign mux_1_61 = (sel[0] == 0)? din122 : din123;
assign mux_1_62 = (sel[0] == 0)? din124 : din125;
assign mux_1_63 = (sel[0] == 0)? din126 : din127;
assign mux_1_64 = (sel[0] == 0)? din128 : din129;
assign mux_1_65 = (sel[0] == 0)? din130 : din131;
assign mux_1_66 = (sel[0] == 0)? din132 : din133;
assign mux_1_67 = (sel[0] == 0)? din134 : din135;
assign mux_1_68 = (sel[0] == 0)? din136 : din137;
assign mux_1_69 = (sel[0] == 0)? din138 : din139;
assign mux_1_70 = (sel[0] == 0)? din140 : din141;
assign mux_1_71 = (sel[0] == 0)? din142 : din143;
assign mux_1_72 = (sel[0] == 0)? din144 : din145;
assign mux_1_73 = (sel[0] == 0)? din146 : din147;
assign mux_1_74 = (sel[0] == 0)? din148 : din149;
assign mux_1_75 = (sel[0] == 0)? din150 : din151;
assign mux_1_76 = (sel[0] == 0)? din152 : din153;
assign mux_1_77 = (sel[0] == 0)? din154 : din155;
assign mux_1_78 = (sel[0] == 0)? din156 : din157;
assign mux_1_79 = (sel[0] == 0)? din158 : din159;
assign mux_1_80 = (sel[0] == 0)? din160 : din161;
assign mux_1_81 = (sel[0] == 0)? din162 : din163;
assign mux_1_82 = (sel[0] == 0)? din164 : din165;
assign mux_1_83 = (sel[0] == 0)? din166 : din167;
assign mux_1_84 = (sel[0] == 0)? din168 : din169;
assign mux_1_85 = (sel[0] == 0)? din170 : din171;
assign mux_1_86 = (sel[0] == 0)? din172 : din173;
assign mux_1_87 = (sel[0] == 0)? din174 : din175;
assign mux_1_88 = (sel[0] == 0)? din176 : din177;
assign mux_1_89 = (sel[0] == 0)? din178 : din179;
assign mux_1_90 = (sel[0] == 0)? din180 : din181;
assign mux_1_91 = (sel[0] == 0)? din182 : din183;
assign mux_1_92 = (sel[0] == 0)? din184 : din185;
assign mux_1_93 = (sel[0] == 0)? din186 : din187;
assign mux_1_94 = (sel[0] == 0)? din188 : din189;
assign mux_1_95 = (sel[0] == 0)? din190 : din191;
assign mux_1_96 = (sel[0] == 0)? din192 : din193;
assign mux_1_97 = (sel[0] == 0)? din194 : din195;
assign mux_1_98 = (sel[0] == 0)? din196 : din197;
assign mux_1_99 = (sel[0] == 0)? din198 : din199;
assign mux_1_100 = (sel[0] == 0)? din200 : din201;
assign mux_1_101 = (sel[0] == 0)? din202 : din203;
assign mux_1_102 = (sel[0] == 0)? din204 : din205;
assign mux_1_103 = (sel[0] == 0)? din206 : din207;
assign mux_1_104 = (sel[0] == 0)? din208 : din209;
assign mux_1_105 = (sel[0] == 0)? din210 : din211;
assign mux_1_106 = (sel[0] == 0)? din212 : din213;
assign mux_1_107 = (sel[0] == 0)? din214 : din215;
assign mux_1_108 = (sel[0] == 0)? din216 : din217;
assign mux_1_109 = (sel[0] == 0)? din218 : din219;
assign mux_1_110 = (sel[0] == 0)? din220 : din221;
assign mux_1_111 = (sel[0] == 0)? din222 : din223;
assign mux_1_112 = (sel[0] == 0)? din224 : din225;
assign mux_1_113 = (sel[0] == 0)? din226 : din227;
assign mux_1_114 = (sel[0] == 0)? din228 : din229;
assign mux_1_115 = (sel[0] == 0)? din230 : din231;
assign mux_1_116 = (sel[0] == 0)? din232 : din233;
assign mux_1_117 = (sel[0] == 0)? din234 : din235;
assign mux_1_118 = (sel[0] == 0)? din236 : din237;
assign mux_1_119 = (sel[0] == 0)? din238 : din239;
assign mux_1_120 = (sel[0] == 0)? din240 : din241;
assign mux_1_121 = (sel[0] == 0)? din242 : din243;
assign mux_1_122 = (sel[0] == 0)? din244 : din245;
assign mux_1_123 = (sel[0] == 0)? din246 : din247;
assign mux_1_124 = (sel[0] == 0)? din248 : din249;
assign mux_1_125 = (sel[0] == 0)? din250 : din251;
assign mux_1_126 = (sel[0] == 0)? din252 : din253;
assign mux_1_127 = (sel[0] == 0)? din254 : din255;
assign mux_1_128 = (sel[0] == 0)? din256 : din257;
assign mux_1_129 = (sel[0] == 0)? din258 : din259;
assign mux_1_130 = (sel[0] == 0)? din260 : din261;
assign mux_1_131 = (sel[0] == 0)? din262 : din263;
assign mux_1_132 = (sel[0] == 0)? din264 : din265;
assign mux_1_133 = (sel[0] == 0)? din266 : din267;
assign mux_1_134 = (sel[0] == 0)? din268 : din269;
assign mux_1_135 = (sel[0] == 0)? din270 : din271;
assign mux_1_136 = (sel[0] == 0)? din272 : din273;
assign mux_1_137 = (sel[0] == 0)? din274 : din275;
assign mux_1_138 = (sel[0] == 0)? din276 : din277;
assign mux_1_139 = (sel[0] == 0)? din278 : din279;
assign mux_1_140 = (sel[0] == 0)? din280 : din281;
assign mux_1_141 = (sel[0] == 0)? din282 : din283;
assign mux_1_142 = (sel[0] == 0)? din284 : din285;
assign mux_1_143 = (sel[0] == 0)? din286 : din287;
assign mux_1_144 = (sel[0] == 0)? din288 : din289;
assign mux_1_145 = (sel[0] == 0)? din290 : din291;
assign mux_1_146 = (sel[0] == 0)? din292 : din293;
assign mux_1_147 = (sel[0] == 0)? din294 : din295;
assign mux_1_148 = (sel[0] == 0)? din296 : din297;
assign mux_1_149 = (sel[0] == 0)? din298 : din299;
assign mux_1_150 = (sel[0] == 0)? din300 : din301;
assign mux_1_151 = (sel[0] == 0)? din302 : din303;
assign mux_1_152 = (sel[0] == 0)? din304 : din305;
assign mux_1_153 = (sel[0] == 0)? din306 : din307;
assign mux_1_154 = (sel[0] == 0)? din308 : din309;
assign mux_1_155 = (sel[0] == 0)? din310 : din311;
assign mux_1_156 = (sel[0] == 0)? din312 : din313;
assign mux_1_157 = (sel[0] == 0)? din314 : din315;
assign mux_1_158 = (sel[0] == 0)? din316 : din317;
assign mux_1_159 = (sel[0] == 0)? din318 : din319;
assign mux_1_160 = (sel[0] == 0)? din320 : din321;
assign mux_1_161 = (sel[0] == 0)? din322 : din323;
assign mux_1_162 = (sel[0] == 0)? din324 : din325;
assign mux_1_163 = (sel[0] == 0)? din326 : din327;
assign mux_1_164 = (sel[0] == 0)? din328 : din329;
assign mux_1_165 = (sel[0] == 0)? din330 : din331;
assign mux_1_166 = (sel[0] == 0)? din332 : din333;
assign mux_1_167 = (sel[0] == 0)? din334 : din335;
assign mux_1_168 = (sel[0] == 0)? din336 : din337;
assign mux_1_169 = (sel[0] == 0)? din338 : din339;
assign mux_1_170 = (sel[0] == 0)? din340 : din341;
assign mux_1_171 = (sel[0] == 0)? din342 : din343;
assign mux_1_172 = (sel[0] == 0)? din344 : din345;
assign mux_1_173 = (sel[0] == 0)? din346 : din347;
assign mux_1_174 = (sel[0] == 0)? din348 : din349;
assign mux_1_175 = (sel[0] == 0)? din350 : din351;
assign mux_1_176 = (sel[0] == 0)? din352 : din353;
assign mux_1_177 = (sel[0] == 0)? din354 : din355;
assign mux_1_178 = (sel[0] == 0)? din356 : din357;
assign mux_1_179 = (sel[0] == 0)? din358 : din359;
assign mux_1_180 = (sel[0] == 0)? din360 : din361;
assign mux_1_181 = (sel[0] == 0)? din362 : din363;
assign mux_1_182 = (sel[0] == 0)? din364 : din365;
assign mux_1_183 = (sel[0] == 0)? din366 : din367;
assign mux_1_184 = (sel[0] == 0)? din368 : din369;
assign mux_1_185 = (sel[0] == 0)? din370 : din371;
assign mux_1_186 = (sel[0] == 0)? din372 : din373;
assign mux_1_187 = (sel[0] == 0)? din374 : din375;
assign mux_1_188 = (sel[0] == 0)? din376 : din377;
assign mux_1_189 = (sel[0] == 0)? din378 : din379;
assign mux_1_190 = (sel[0] == 0)? din380 : din381;
assign mux_1_191 = (sel[0] == 0)? din382 : din383;
assign mux_1_192 = (sel[0] == 0)? din384 : din385;
assign mux_1_193 = (sel[0] == 0)? din386 : din387;
assign mux_1_194 = (sel[0] == 0)? din388 : din389;
assign mux_1_195 = (sel[0] == 0)? din390 : din391;
assign mux_1_196 = (sel[0] == 0)? din392 : din393;
assign mux_1_197 = (sel[0] == 0)? din394 : din395;
assign mux_1_198 = (sel[0] == 0)? din396 : din397;
assign mux_1_199 = (sel[0] == 0)? din398 : din399;
assign mux_1_200 = (sel[0] == 0)? din400 : din401;
assign mux_1_201 = (sel[0] == 0)? din402 : din403;
assign mux_1_202 = (sel[0] == 0)? din404 : din405;
assign mux_1_203 = (sel[0] == 0)? din406 : din407;
assign mux_1_204 = (sel[0] == 0)? din408 : din409;
assign mux_1_205 = (sel[0] == 0)? din410 : din411;
assign mux_1_206 = (sel[0] == 0)? din412 : din413;
assign mux_1_207 = (sel[0] == 0)? din414 : din415;
assign mux_1_208 = (sel[0] == 0)? din416 : din417;
assign mux_1_209 = (sel[0] == 0)? din418 : din419;
assign mux_1_210 = (sel[0] == 0)? din420 : din421;
assign mux_1_211 = (sel[0] == 0)? din422 : din423;
assign mux_1_212 = (sel[0] == 0)? din424 : din425;
assign mux_1_213 = (sel[0] == 0)? din426 : din427;
assign mux_1_214 = (sel[0] == 0)? din428 : din429;
assign mux_1_215 = (sel[0] == 0)? din430 : din431;
assign mux_1_216 = (sel[0] == 0)? din432 : din433;
assign mux_1_217 = (sel[0] == 0)? din434 : din435;
assign mux_1_218 = (sel[0] == 0)? din436 : din437;
assign mux_1_219 = (sel[0] == 0)? din438 : din439;
assign mux_1_220 = (sel[0] == 0)? din440 : din441;
assign mux_1_221 = (sel[0] == 0)? din442 : din443;
assign mux_1_222 = (sel[0] == 0)? din444 : din445;
assign mux_1_223 = (sel[0] == 0)? din446 : din447;
assign mux_1_224 = (sel[0] == 0)? din448 : din449;
assign mux_1_225 = (sel[0] == 0)? din450 : din451;
assign mux_1_226 = (sel[0] == 0)? din452 : din453;
assign mux_1_227 = (sel[0] == 0)? din454 : din455;
assign mux_1_228 = (sel[0] == 0)? din456 : din457;
assign mux_1_229 = (sel[0] == 0)? din458 : din459;
assign mux_1_230 = (sel[0] == 0)? din460 : din461;
assign mux_1_231 = (sel[0] == 0)? din462 : din463;
assign mux_1_232 = (sel[0] == 0)? din464 : din465;
assign mux_1_233 = (sel[0] == 0)? din466 : din467;
assign mux_1_234 = (sel[0] == 0)? din468 : din469;
assign mux_1_235 = (sel[0] == 0)? din470 : din471;
assign mux_1_236 = (sel[0] == 0)? din472 : din473;
assign mux_1_237 = (sel[0] == 0)? din474 : din475;
assign mux_1_238 = (sel[0] == 0)? din476 : din477;
assign mux_1_239 = (sel[0] == 0)? din478 : din479;
assign mux_1_240 = (sel[0] == 0)? din480 : din481;
assign mux_1_241 = (sel[0] == 0)? din482 : din483;
assign mux_1_242 = (sel[0] == 0)? din484 : din485;
assign mux_1_243 = (sel[0] == 0)? din486 : din487;
assign mux_1_244 = (sel[0] == 0)? din488 : din489;
assign mux_1_245 = (sel[0] == 0)? din490 : din491;
assign mux_1_246 = (sel[0] == 0)? din492 : din493;
assign mux_1_247 = (sel[0] == 0)? din494 : din495;
assign mux_1_248 = (sel[0] == 0)? din496 : din497;
assign mux_1_249 = (sel[0] == 0)? din498 : din499;
assign mux_1_250 = (sel[0] == 0)? din500 : din501;
assign mux_1_251 = (sel[0] == 0)? din502 : din503;
assign mux_1_252 = (sel[0] == 0)? din504 : din505;
assign mux_1_253 = (sel[0] == 0)? din506 : din507;
assign mux_1_254 = (sel[0] == 0)? din508 : din509;
assign mux_1_255 = (sel[0] == 0)? din510 : din511;
assign mux_1_256 = (sel[0] == 0)? din512 : din513;
assign mux_1_257 = (sel[0] == 0)? din514 : din515;
assign mux_1_258 = (sel[0] == 0)? din516 : din517;
assign mux_1_259 = (sel[0] == 0)? din518 : din519;
assign mux_1_260 = (sel[0] == 0)? din520 : din521;
assign mux_1_261 = (sel[0] == 0)? din522 : din523;
assign mux_1_262 = (sel[0] == 0)? din524 : din525;
assign mux_1_263 = (sel[0] == 0)? din526 : din527;
assign mux_1_264 = (sel[0] == 0)? din528 : din529;
assign mux_1_265 = (sel[0] == 0)? din530 : din531;
assign mux_1_266 = (sel[0] == 0)? din532 : din533;
assign mux_1_267 = (sel[0] == 0)? din534 : din535;
assign mux_1_268 = (sel[0] == 0)? din536 : din537;
assign mux_1_269 = (sel[0] == 0)? din538 : din539;
assign mux_1_270 = (sel[0] == 0)? din540 : din541;
assign mux_1_271 = (sel[0] == 0)? din542 : din543;
assign mux_1_272 = (sel[0] == 0)? din544 : din545;
assign mux_1_273 = (sel[0] == 0)? din546 : din547;
assign mux_1_274 = (sel[0] == 0)? din548 : din549;
assign mux_1_275 = (sel[0] == 0)? din550 : din551;
assign mux_1_276 = (sel[0] == 0)? din552 : din553;
assign mux_1_277 = (sel[0] == 0)? din554 : din555;
assign mux_1_278 = (sel[0] == 0)? din556 : din557;
assign mux_1_279 = (sel[0] == 0)? din558 : din559;
assign mux_1_280 = (sel[0] == 0)? din560 : din561;
assign mux_1_281 = (sel[0] == 0)? din562 : din563;
assign mux_1_282 = (sel[0] == 0)? din564 : din565;
assign mux_1_283 = (sel[0] == 0)? din566 : din567;
assign mux_1_284 = (sel[0] == 0)? din568 : din569;
assign mux_1_285 = (sel[0] == 0)? din570 : din571;
assign mux_1_286 = (sel[0] == 0)? din572 : din573;
assign mux_1_287 = (sel[0] == 0)? din574 : din575;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;
assign mux_2_1 = (sel[1] == 0)? mux_1_2 : mux_1_3;
assign mux_2_2 = (sel[1] == 0)? mux_1_4 : mux_1_5;
assign mux_2_3 = (sel[1] == 0)? mux_1_6 : mux_1_7;
assign mux_2_4 = (sel[1] == 0)? mux_1_8 : mux_1_9;
assign mux_2_5 = (sel[1] == 0)? mux_1_10 : mux_1_11;
assign mux_2_6 = (sel[1] == 0)? mux_1_12 : mux_1_13;
assign mux_2_7 = (sel[1] == 0)? mux_1_14 : mux_1_15;
assign mux_2_8 = (sel[1] == 0)? mux_1_16 : mux_1_17;
assign mux_2_9 = (sel[1] == 0)? mux_1_18 : mux_1_19;
assign mux_2_10 = (sel[1] == 0)? mux_1_20 : mux_1_21;
assign mux_2_11 = (sel[1] == 0)? mux_1_22 : mux_1_23;
assign mux_2_12 = (sel[1] == 0)? mux_1_24 : mux_1_25;
assign mux_2_13 = (sel[1] == 0)? mux_1_26 : mux_1_27;
assign mux_2_14 = (sel[1] == 0)? mux_1_28 : mux_1_29;
assign mux_2_15 = (sel[1] == 0)? mux_1_30 : mux_1_31;
assign mux_2_16 = (sel[1] == 0)? mux_1_32 : mux_1_33;
assign mux_2_17 = (sel[1] == 0)? mux_1_34 : mux_1_35;
assign mux_2_18 = (sel[1] == 0)? mux_1_36 : mux_1_37;
assign mux_2_19 = (sel[1] == 0)? mux_1_38 : mux_1_39;
assign mux_2_20 = (sel[1] == 0)? mux_1_40 : mux_1_41;
assign mux_2_21 = (sel[1] == 0)? mux_1_42 : mux_1_43;
assign mux_2_22 = (sel[1] == 0)? mux_1_44 : mux_1_45;
assign mux_2_23 = (sel[1] == 0)? mux_1_46 : mux_1_47;
assign mux_2_24 = (sel[1] == 0)? mux_1_48 : mux_1_49;
assign mux_2_25 = (sel[1] == 0)? mux_1_50 : mux_1_51;
assign mux_2_26 = (sel[1] == 0)? mux_1_52 : mux_1_53;
assign mux_2_27 = (sel[1] == 0)? mux_1_54 : mux_1_55;
assign mux_2_28 = (sel[1] == 0)? mux_1_56 : mux_1_57;
assign mux_2_29 = (sel[1] == 0)? mux_1_58 : mux_1_59;
assign mux_2_30 = (sel[1] == 0)? mux_1_60 : mux_1_61;
assign mux_2_31 = (sel[1] == 0)? mux_1_62 : mux_1_63;
assign mux_2_32 = (sel[1] == 0)? mux_1_64 : mux_1_65;
assign mux_2_33 = (sel[1] == 0)? mux_1_66 : mux_1_67;
assign mux_2_34 = (sel[1] == 0)? mux_1_68 : mux_1_69;
assign mux_2_35 = (sel[1] == 0)? mux_1_70 : mux_1_71;
assign mux_2_36 = (sel[1] == 0)? mux_1_72 : mux_1_73;
assign mux_2_37 = (sel[1] == 0)? mux_1_74 : mux_1_75;
assign mux_2_38 = (sel[1] == 0)? mux_1_76 : mux_1_77;
assign mux_2_39 = (sel[1] == 0)? mux_1_78 : mux_1_79;
assign mux_2_40 = (sel[1] == 0)? mux_1_80 : mux_1_81;
assign mux_2_41 = (sel[1] == 0)? mux_1_82 : mux_1_83;
assign mux_2_42 = (sel[1] == 0)? mux_1_84 : mux_1_85;
assign mux_2_43 = (sel[1] == 0)? mux_1_86 : mux_1_87;
assign mux_2_44 = (sel[1] == 0)? mux_1_88 : mux_1_89;
assign mux_2_45 = (sel[1] == 0)? mux_1_90 : mux_1_91;
assign mux_2_46 = (sel[1] == 0)? mux_1_92 : mux_1_93;
assign mux_2_47 = (sel[1] == 0)? mux_1_94 : mux_1_95;
assign mux_2_48 = (sel[1] == 0)? mux_1_96 : mux_1_97;
assign mux_2_49 = (sel[1] == 0)? mux_1_98 : mux_1_99;
assign mux_2_50 = (sel[1] == 0)? mux_1_100 : mux_1_101;
assign mux_2_51 = (sel[1] == 0)? mux_1_102 : mux_1_103;
assign mux_2_52 = (sel[1] == 0)? mux_1_104 : mux_1_105;
assign mux_2_53 = (sel[1] == 0)? mux_1_106 : mux_1_107;
assign mux_2_54 = (sel[1] == 0)? mux_1_108 : mux_1_109;
assign mux_2_55 = (sel[1] == 0)? mux_1_110 : mux_1_111;
assign mux_2_56 = (sel[1] == 0)? mux_1_112 : mux_1_113;
assign mux_2_57 = (sel[1] == 0)? mux_1_114 : mux_1_115;
assign mux_2_58 = (sel[1] == 0)? mux_1_116 : mux_1_117;
assign mux_2_59 = (sel[1] == 0)? mux_1_118 : mux_1_119;
assign mux_2_60 = (sel[1] == 0)? mux_1_120 : mux_1_121;
assign mux_2_61 = (sel[1] == 0)? mux_1_122 : mux_1_123;
assign mux_2_62 = (sel[1] == 0)? mux_1_124 : mux_1_125;
assign mux_2_63 = (sel[1] == 0)? mux_1_126 : mux_1_127;
assign mux_2_64 = (sel[1] == 0)? mux_1_128 : mux_1_129;
assign mux_2_65 = (sel[1] == 0)? mux_1_130 : mux_1_131;
assign mux_2_66 = (sel[1] == 0)? mux_1_132 : mux_1_133;
assign mux_2_67 = (sel[1] == 0)? mux_1_134 : mux_1_135;
assign mux_2_68 = (sel[1] == 0)? mux_1_136 : mux_1_137;
assign mux_2_69 = (sel[1] == 0)? mux_1_138 : mux_1_139;
assign mux_2_70 = (sel[1] == 0)? mux_1_140 : mux_1_141;
assign mux_2_71 = (sel[1] == 0)? mux_1_142 : mux_1_143;
assign mux_2_72 = (sel[1] == 0)? mux_1_144 : mux_1_145;
assign mux_2_73 = (sel[1] == 0)? mux_1_146 : mux_1_147;
assign mux_2_74 = (sel[1] == 0)? mux_1_148 : mux_1_149;
assign mux_2_75 = (sel[1] == 0)? mux_1_150 : mux_1_151;
assign mux_2_76 = (sel[1] == 0)? mux_1_152 : mux_1_153;
assign mux_2_77 = (sel[1] == 0)? mux_1_154 : mux_1_155;
assign mux_2_78 = (sel[1] == 0)? mux_1_156 : mux_1_157;
assign mux_2_79 = (sel[1] == 0)? mux_1_158 : mux_1_159;
assign mux_2_80 = (sel[1] == 0)? mux_1_160 : mux_1_161;
assign mux_2_81 = (sel[1] == 0)? mux_1_162 : mux_1_163;
assign mux_2_82 = (sel[1] == 0)? mux_1_164 : mux_1_165;
assign mux_2_83 = (sel[1] == 0)? mux_1_166 : mux_1_167;
assign mux_2_84 = (sel[1] == 0)? mux_1_168 : mux_1_169;
assign mux_2_85 = (sel[1] == 0)? mux_1_170 : mux_1_171;
assign mux_2_86 = (sel[1] == 0)? mux_1_172 : mux_1_173;
assign mux_2_87 = (sel[1] == 0)? mux_1_174 : mux_1_175;
assign mux_2_88 = (sel[1] == 0)? mux_1_176 : mux_1_177;
assign mux_2_89 = (sel[1] == 0)? mux_1_178 : mux_1_179;
assign mux_2_90 = (sel[1] == 0)? mux_1_180 : mux_1_181;
assign mux_2_91 = (sel[1] == 0)? mux_1_182 : mux_1_183;
assign mux_2_92 = (sel[1] == 0)? mux_1_184 : mux_1_185;
assign mux_2_93 = (sel[1] == 0)? mux_1_186 : mux_1_187;
assign mux_2_94 = (sel[1] == 0)? mux_1_188 : mux_1_189;
assign mux_2_95 = (sel[1] == 0)? mux_1_190 : mux_1_191;
assign mux_2_96 = (sel[1] == 0)? mux_1_192 : mux_1_193;
assign mux_2_97 = (sel[1] == 0)? mux_1_194 : mux_1_195;
assign mux_2_98 = (sel[1] == 0)? mux_1_196 : mux_1_197;
assign mux_2_99 = (sel[1] == 0)? mux_1_198 : mux_1_199;
assign mux_2_100 = (sel[1] == 0)? mux_1_200 : mux_1_201;
assign mux_2_101 = (sel[1] == 0)? mux_1_202 : mux_1_203;
assign mux_2_102 = (sel[1] == 0)? mux_1_204 : mux_1_205;
assign mux_2_103 = (sel[1] == 0)? mux_1_206 : mux_1_207;
assign mux_2_104 = (sel[1] == 0)? mux_1_208 : mux_1_209;
assign mux_2_105 = (sel[1] == 0)? mux_1_210 : mux_1_211;
assign mux_2_106 = (sel[1] == 0)? mux_1_212 : mux_1_213;
assign mux_2_107 = (sel[1] == 0)? mux_1_214 : mux_1_215;
assign mux_2_108 = (sel[1] == 0)? mux_1_216 : mux_1_217;
assign mux_2_109 = (sel[1] == 0)? mux_1_218 : mux_1_219;
assign mux_2_110 = (sel[1] == 0)? mux_1_220 : mux_1_221;
assign mux_2_111 = (sel[1] == 0)? mux_1_222 : mux_1_223;
assign mux_2_112 = (sel[1] == 0)? mux_1_224 : mux_1_225;
assign mux_2_113 = (sel[1] == 0)? mux_1_226 : mux_1_227;
assign mux_2_114 = (sel[1] == 0)? mux_1_228 : mux_1_229;
assign mux_2_115 = (sel[1] == 0)? mux_1_230 : mux_1_231;
assign mux_2_116 = (sel[1] == 0)? mux_1_232 : mux_1_233;
assign mux_2_117 = (sel[1] == 0)? mux_1_234 : mux_1_235;
assign mux_2_118 = (sel[1] == 0)? mux_1_236 : mux_1_237;
assign mux_2_119 = (sel[1] == 0)? mux_1_238 : mux_1_239;
assign mux_2_120 = (sel[1] == 0)? mux_1_240 : mux_1_241;
assign mux_2_121 = (sel[1] == 0)? mux_1_242 : mux_1_243;
assign mux_2_122 = (sel[1] == 0)? mux_1_244 : mux_1_245;
assign mux_2_123 = (sel[1] == 0)? mux_1_246 : mux_1_247;
assign mux_2_124 = (sel[1] == 0)? mux_1_248 : mux_1_249;
assign mux_2_125 = (sel[1] == 0)? mux_1_250 : mux_1_251;
assign mux_2_126 = (sel[1] == 0)? mux_1_252 : mux_1_253;
assign mux_2_127 = (sel[1] == 0)? mux_1_254 : mux_1_255;
assign mux_2_128 = (sel[1] == 0)? mux_1_256 : mux_1_257;
assign mux_2_129 = (sel[1] == 0)? mux_1_258 : mux_1_259;
assign mux_2_130 = (sel[1] == 0)? mux_1_260 : mux_1_261;
assign mux_2_131 = (sel[1] == 0)? mux_1_262 : mux_1_263;
assign mux_2_132 = (sel[1] == 0)? mux_1_264 : mux_1_265;
assign mux_2_133 = (sel[1] == 0)? mux_1_266 : mux_1_267;
assign mux_2_134 = (sel[1] == 0)? mux_1_268 : mux_1_269;
assign mux_2_135 = (sel[1] == 0)? mux_1_270 : mux_1_271;
assign mux_2_136 = (sel[1] == 0)? mux_1_272 : mux_1_273;
assign mux_2_137 = (sel[1] == 0)? mux_1_274 : mux_1_275;
assign mux_2_138 = (sel[1] == 0)? mux_1_276 : mux_1_277;
assign mux_2_139 = (sel[1] == 0)? mux_1_278 : mux_1_279;
assign mux_2_140 = (sel[1] == 0)? mux_1_280 : mux_1_281;
assign mux_2_141 = (sel[1] == 0)? mux_1_282 : mux_1_283;
assign mux_2_142 = (sel[1] == 0)? mux_1_284 : mux_1_285;
assign mux_2_143 = (sel[1] == 0)? mux_1_286 : mux_1_287;

// Generate level 3 logic
assign mux_3_0 = (sel[2] == 0)? mux_2_0 : mux_2_1;
assign mux_3_1 = (sel[2] == 0)? mux_2_2 : mux_2_3;
assign mux_3_2 = (sel[2] == 0)? mux_2_4 : mux_2_5;
assign mux_3_3 = (sel[2] == 0)? mux_2_6 : mux_2_7;
assign mux_3_4 = (sel[2] == 0)? mux_2_8 : mux_2_9;
assign mux_3_5 = (sel[2] == 0)? mux_2_10 : mux_2_11;
assign mux_3_6 = (sel[2] == 0)? mux_2_12 : mux_2_13;
assign mux_3_7 = (sel[2] == 0)? mux_2_14 : mux_2_15;
assign mux_3_8 = (sel[2] == 0)? mux_2_16 : mux_2_17;
assign mux_3_9 = (sel[2] == 0)? mux_2_18 : mux_2_19;
assign mux_3_10 = (sel[2] == 0)? mux_2_20 : mux_2_21;
assign mux_3_11 = (sel[2] == 0)? mux_2_22 : mux_2_23;
assign mux_3_12 = (sel[2] == 0)? mux_2_24 : mux_2_25;
assign mux_3_13 = (sel[2] == 0)? mux_2_26 : mux_2_27;
assign mux_3_14 = (sel[2] == 0)? mux_2_28 : mux_2_29;
assign mux_3_15 = (sel[2] == 0)? mux_2_30 : mux_2_31;
assign mux_3_16 = (sel[2] == 0)? mux_2_32 : mux_2_33;
assign mux_3_17 = (sel[2] == 0)? mux_2_34 : mux_2_35;
assign mux_3_18 = (sel[2] == 0)? mux_2_36 : mux_2_37;
assign mux_3_19 = (sel[2] == 0)? mux_2_38 : mux_2_39;
assign mux_3_20 = (sel[2] == 0)? mux_2_40 : mux_2_41;
assign mux_3_21 = (sel[2] == 0)? mux_2_42 : mux_2_43;
assign mux_3_22 = (sel[2] == 0)? mux_2_44 : mux_2_45;
assign mux_3_23 = (sel[2] == 0)? mux_2_46 : mux_2_47;
assign mux_3_24 = (sel[2] == 0)? mux_2_48 : mux_2_49;
assign mux_3_25 = (sel[2] == 0)? mux_2_50 : mux_2_51;
assign mux_3_26 = (sel[2] == 0)? mux_2_52 : mux_2_53;
assign mux_3_27 = (sel[2] == 0)? mux_2_54 : mux_2_55;
assign mux_3_28 = (sel[2] == 0)? mux_2_56 : mux_2_57;
assign mux_3_29 = (sel[2] == 0)? mux_2_58 : mux_2_59;
assign mux_3_30 = (sel[2] == 0)? mux_2_60 : mux_2_61;
assign mux_3_31 = (sel[2] == 0)? mux_2_62 : mux_2_63;
assign mux_3_32 = (sel[2] == 0)? mux_2_64 : mux_2_65;
assign mux_3_33 = (sel[2] == 0)? mux_2_66 : mux_2_67;
assign mux_3_34 = (sel[2] == 0)? mux_2_68 : mux_2_69;
assign mux_3_35 = (sel[2] == 0)? mux_2_70 : mux_2_71;
assign mux_3_36 = (sel[2] == 0)? mux_2_72 : mux_2_73;
assign mux_3_37 = (sel[2] == 0)? mux_2_74 : mux_2_75;
assign mux_3_38 = (sel[2] == 0)? mux_2_76 : mux_2_77;
assign mux_3_39 = (sel[2] == 0)? mux_2_78 : mux_2_79;
assign mux_3_40 = (sel[2] == 0)? mux_2_80 : mux_2_81;
assign mux_3_41 = (sel[2] == 0)? mux_2_82 : mux_2_83;
assign mux_3_42 = (sel[2] == 0)? mux_2_84 : mux_2_85;
assign mux_3_43 = (sel[2] == 0)? mux_2_86 : mux_2_87;
assign mux_3_44 = (sel[2] == 0)? mux_2_88 : mux_2_89;
assign mux_3_45 = (sel[2] == 0)? mux_2_90 : mux_2_91;
assign mux_3_46 = (sel[2] == 0)? mux_2_92 : mux_2_93;
assign mux_3_47 = (sel[2] == 0)? mux_2_94 : mux_2_95;
assign mux_3_48 = (sel[2] == 0)? mux_2_96 : mux_2_97;
assign mux_3_49 = (sel[2] == 0)? mux_2_98 : mux_2_99;
assign mux_3_50 = (sel[2] == 0)? mux_2_100 : mux_2_101;
assign mux_3_51 = (sel[2] == 0)? mux_2_102 : mux_2_103;
assign mux_3_52 = (sel[2] == 0)? mux_2_104 : mux_2_105;
assign mux_3_53 = (sel[2] == 0)? mux_2_106 : mux_2_107;
assign mux_3_54 = (sel[2] == 0)? mux_2_108 : mux_2_109;
assign mux_3_55 = (sel[2] == 0)? mux_2_110 : mux_2_111;
assign mux_3_56 = (sel[2] == 0)? mux_2_112 : mux_2_113;
assign mux_3_57 = (sel[2] == 0)? mux_2_114 : mux_2_115;
assign mux_3_58 = (sel[2] == 0)? mux_2_116 : mux_2_117;
assign mux_3_59 = (sel[2] == 0)? mux_2_118 : mux_2_119;
assign mux_3_60 = (sel[2] == 0)? mux_2_120 : mux_2_121;
assign mux_3_61 = (sel[2] == 0)? mux_2_122 : mux_2_123;
assign mux_3_62 = (sel[2] == 0)? mux_2_124 : mux_2_125;
assign mux_3_63 = (sel[2] == 0)? mux_2_126 : mux_2_127;
assign mux_3_64 = (sel[2] == 0)? mux_2_128 : mux_2_129;
assign mux_3_65 = (sel[2] == 0)? mux_2_130 : mux_2_131;
assign mux_3_66 = (sel[2] == 0)? mux_2_132 : mux_2_133;
assign mux_3_67 = (sel[2] == 0)? mux_2_134 : mux_2_135;
assign mux_3_68 = (sel[2] == 0)? mux_2_136 : mux_2_137;
assign mux_3_69 = (sel[2] == 0)? mux_2_138 : mux_2_139;
assign mux_3_70 = (sel[2] == 0)? mux_2_140 : mux_2_141;
assign mux_3_71 = (sel[2] == 0)? mux_2_142 : mux_2_143;

// Generate level 4 logic
assign mux_4_0 = (sel[3] == 0)? mux_3_0 : mux_3_1;
assign mux_4_1 = (sel[3] == 0)? mux_3_2 : mux_3_3;
assign mux_4_2 = (sel[3] == 0)? mux_3_4 : mux_3_5;
assign mux_4_3 = (sel[3] == 0)? mux_3_6 : mux_3_7;
assign mux_4_4 = (sel[3] == 0)? mux_3_8 : mux_3_9;
assign mux_4_5 = (sel[3] == 0)? mux_3_10 : mux_3_11;
assign mux_4_6 = (sel[3] == 0)? mux_3_12 : mux_3_13;
assign mux_4_7 = (sel[3] == 0)? mux_3_14 : mux_3_15;
assign mux_4_8 = (sel[3] == 0)? mux_3_16 : mux_3_17;
assign mux_4_9 = (sel[3] == 0)? mux_3_18 : mux_3_19;
assign mux_4_10 = (sel[3] == 0)? mux_3_20 : mux_3_21;
assign mux_4_11 = (sel[3] == 0)? mux_3_22 : mux_3_23;
assign mux_4_12 = (sel[3] == 0)? mux_3_24 : mux_3_25;
assign mux_4_13 = (sel[3] == 0)? mux_3_26 : mux_3_27;
assign mux_4_14 = (sel[3] == 0)? mux_3_28 : mux_3_29;
assign mux_4_15 = (sel[3] == 0)? mux_3_30 : mux_3_31;
assign mux_4_16 = (sel[3] == 0)? mux_3_32 : mux_3_33;
assign mux_4_17 = (sel[3] == 0)? mux_3_34 : mux_3_35;
assign mux_4_18 = (sel[3] == 0)? mux_3_36 : mux_3_37;
assign mux_4_19 = (sel[3] == 0)? mux_3_38 : mux_3_39;
assign mux_4_20 = (sel[3] == 0)? mux_3_40 : mux_3_41;
assign mux_4_21 = (sel[3] == 0)? mux_3_42 : mux_3_43;
assign mux_4_22 = (sel[3] == 0)? mux_3_44 : mux_3_45;
assign mux_4_23 = (sel[3] == 0)? mux_3_46 : mux_3_47;
assign mux_4_24 = (sel[3] == 0)? mux_3_48 : mux_3_49;
assign mux_4_25 = (sel[3] == 0)? mux_3_50 : mux_3_51;
assign mux_4_26 = (sel[3] == 0)? mux_3_52 : mux_3_53;
assign mux_4_27 = (sel[3] == 0)? mux_3_54 : mux_3_55;
assign mux_4_28 = (sel[3] == 0)? mux_3_56 : mux_3_57;
assign mux_4_29 = (sel[3] == 0)? mux_3_58 : mux_3_59;
assign mux_4_30 = (sel[3] == 0)? mux_3_60 : mux_3_61;
assign mux_4_31 = (sel[3] == 0)? mux_3_62 : mux_3_63;
assign mux_4_32 = (sel[3] == 0)? mux_3_64 : mux_3_65;
assign mux_4_33 = (sel[3] == 0)? mux_3_66 : mux_3_67;
assign mux_4_34 = (sel[3] == 0)? mux_3_68 : mux_3_69;
assign mux_4_35 = (sel[3] == 0)? mux_3_70 : mux_3_71;

// Generate level 5 logic
assign mux_5_0 = (sel[4] == 0)? mux_4_0 : mux_4_1;
assign mux_5_1 = (sel[4] == 0)? mux_4_2 : mux_4_3;
assign mux_5_2 = (sel[4] == 0)? mux_4_4 : mux_4_5;
assign mux_5_3 = (sel[4] == 0)? mux_4_6 : mux_4_7;
assign mux_5_4 = (sel[4] == 0)? mux_4_8 : mux_4_9;
assign mux_5_5 = (sel[4] == 0)? mux_4_10 : mux_4_11;
assign mux_5_6 = (sel[4] == 0)? mux_4_12 : mux_4_13;
assign mux_5_7 = (sel[4] == 0)? mux_4_14 : mux_4_15;
assign mux_5_8 = (sel[4] == 0)? mux_4_16 : mux_4_17;
assign mux_5_9 = (sel[4] == 0)? mux_4_18 : mux_4_19;
assign mux_5_10 = (sel[4] == 0)? mux_4_20 : mux_4_21;
assign mux_5_11 = (sel[4] == 0)? mux_4_22 : mux_4_23;
assign mux_5_12 = (sel[4] == 0)? mux_4_24 : mux_4_25;
assign mux_5_13 = (sel[4] == 0)? mux_4_26 : mux_4_27;
assign mux_5_14 = (sel[4] == 0)? mux_4_28 : mux_4_29;
assign mux_5_15 = (sel[4] == 0)? mux_4_30 : mux_4_31;
assign mux_5_16 = (sel[4] == 0)? mux_4_32 : mux_4_33;
assign mux_5_17 = (sel[4] == 0)? mux_4_34 : mux_4_35;

// Generate level 6 logic
assign mux_6_0 = (sel[5] == 0)? mux_5_0 : mux_5_1;
assign mux_6_1 = (sel[5] == 0)? mux_5_2 : mux_5_3;
assign mux_6_2 = (sel[5] == 0)? mux_5_4 : mux_5_5;
assign mux_6_3 = (sel[5] == 0)? mux_5_6 : mux_5_7;
assign mux_6_4 = (sel[5] == 0)? mux_5_8 : mux_5_9;
assign mux_6_5 = (sel[5] == 0)? mux_5_10 : mux_5_11;
assign mux_6_6 = (sel[5] == 0)? mux_5_12 : mux_5_13;
assign mux_6_7 = (sel[5] == 0)? mux_5_14 : mux_5_15;
assign mux_6_8 = (sel[5] == 0)? mux_5_16 : mux_5_17;

// Generate level 7 logic
assign mux_7_0 = (sel[6] == 0)? mux_6_0 : mux_6_1;
assign mux_7_1 = (sel[6] == 0)? mux_6_2 : mux_6_3;
assign mux_7_2 = (sel[6] == 0)? mux_6_4 : mux_6_5;
assign mux_7_3 = (sel[6] == 0)? mux_6_6 : mux_6_7;
assign mux_7_4 = mux_6_8;

// Generate level 8 logic
assign mux_8_0 = (sel[7] == 0)? mux_7_0 : mux_7_1;
assign mux_8_1 = (sel[7] == 0)? mux_7_2 : mux_7_3;
assign mux_8_2 = mux_7_4;

// Generate level 9 logic
assign mux_9_0 = (sel[8] == 0)? mux_8_0 : mux_8_1;
assign mux_9_1 = mux_8_2;

// Generate level 10 logic
assign mux_10_0 = (sel[9] == 0)? mux_9_0 : mux_9_1;

// output logic
assign dout = mux_10_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActdEe.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActdEe_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActdEe_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActdEe(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActdEe_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActdEe_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdbE.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcdbE_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdbE_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcdbE(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcdbE_rom Thresholding_Batch_0_Thresholding_BatcdbE_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccRA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccRA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccRA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccRA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccRA_rom Thresholding_Batch_0_Thresholding_BatccRA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccVB.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccVB_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccVB_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccVB(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccVB_rom Thresholding_Batch_0_Thresholding_BatccVB_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbtn.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbtn_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbtn_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbtn(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbtn_rom Thresholding_Batch_0_Thresholding_Batcbtn_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/209a/hdl/ramb18_sdp.v

/*
 Copyright (c) 2020, Xilinx
 All rights reserved.

 Redistribution and use in source and binary forms, with or without
 modification, are permitted provided that the following conditions are met:

 * Redistributions of source code must retain the above copyright notice, this
   list of conditions and the following disclaimer.

 * Redistributions in binary form must reproduce the above copyright notice,
   this list of conditions and the following disclaimer in the documentation
   and/or other materials provided with the distribution.

 * Neither the name of FINN nor the names of its
   contributors may be used to endorse or promote products derived from
   this software without specific prior written permission.

 THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
 FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
 SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
 CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
 OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

module ramb18_sdp
#(
    parameter ID = 0,
    parameter DWIDTH = 18,
    parameter AWIDTH = 10,
    parameter DEPTH = 2**AWIDTH,
    parameter MEM_INIT = "",
    parameter RAM_STYLE = "auto"
)
(
	input clk,

	input ena,
	input wea,
	input [AWIDTH-1:0] addra,
	input [DWIDTH-1:0] wdataa,

    input enb,
    input enqb,
	input [AWIDTH-1:0] addrb,
	output reg [DWIDTH-1:0] rdqb
);

(* ram_style = RAM_STYLE *) reg [DWIDTH-1:0] mem[0:DEPTH-1];
reg [DWIDTH-1:0] rdatab;

`ifdef SYNTHESIS
reg [7:0] idx = ID;
`else
reg [15:0] idx;
`endif

//initialize memory
initial begin
  //note the hacky way of adding a filename memblock_ID.dat to the path provided in MEM_INIT
  //ID can go up to 99
  if (ID < 0 && ID > 99) begin
    $display("ID out of range [0-99]");
    $finish();
  end
	//MEM_INIT path must be terminated by /
  `ifdef SYNTHESIS
  if (ID < 10)
    $readmemh({MEM_INIT,"memblock_",idx+8'd48,".dat"}, mem, 0, DEPTH-1);
  else
    $readmemh({MEM_INIT,"memblock_",(idx/10)+8'd48,(idx%10)+8'd48,".dat"}, mem, 0, DEPTH-1);
  `else
  $sformat(idx,"%0d",ID);
  if (ID < 10)
    $readmemh({MEM_INIT,"memblock_",idx[7:0],".dat"}, mem, 0, DEPTH-1);
  else
    $readmemh({MEM_INIT,"memblock_",idx,".dat"}, mem, 0, DEPTH-1);
  `endif
end

//memory ports, with output pipeline register
always @(posedge clk) begin
    if(wea)
        mem[addra] <= wdataa;
    if(enb)
        rdatab <= mem[addrb];
    if(enqb)
        rdqb <= rdatab;
end

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActjbC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActjbC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActjbC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActjbC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActjbC_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActjbC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcddE.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcddE_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcddE_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcddE(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcddE_rom Thresholding_Batch_0_Thresholding_BatcddE_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc9D.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcc9D_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc9D_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcc9D(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcc9D_rom Thresholding_Batch_0_Thresholding_Batcc9D_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/5609/StreamingFIFO_1.v


module StreamingFIFO_1(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [7:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(8)
)
StreamingFIFO_1_StreamingFIFO_1
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActMgi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActMgi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActMgi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActMgi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActMgi_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActMgi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcciv.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcciv_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcciv_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcciv(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcciv_rom Thresholding_Batch_0_Thresholding_Batcciv_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActqcK.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActqcK_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActqcK_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActqcK(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActqcK_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActqcK_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActQgW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActQgW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActQgW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActQgW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActQgW_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActQgW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccTB.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccTB_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccTB_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccTB(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccTB_rom Thresholding_Batch_0_Thresholding_BatccTB_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actbkb_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actbkb_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actbkb(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actbkb_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actbkb_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActGfk.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActGfk_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActGfk_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActGfk(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActGfk_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActGfk_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcrcU.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcrcU_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 5;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcrcU_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcrcU(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd5;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcrcU_rom Thresholding_Batch_0_Thresholding_BatcrcU_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Act2iS.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Act2iS_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Act2iS_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Act2iS(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Act2iS_rom StreamingFCLayer_Batch_4_Matrix_Vector_Act2iS_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Acttde.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Acttde_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Acttde_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Acttde(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Acttde_rom StreamingFCLayer_Batch_1_Matrix_Vector_Acttde_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Act3i2.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Act3i2_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Act3i2_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Act3i2(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Act3i2_rom StreamingFCLayer_Batch_4_Matrix_Vector_Act3i2_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActIfE.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActIfE_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActIfE_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActIfE(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActIfE_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActIfE_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccUB.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccUB_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccUB_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccUB(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccUB_rom Thresholding_Batch_0_Thresholding_BatccUB_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8b1e/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc5D.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcc5D_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc5D_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcc5D(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcc5D_rom Thresholding_Batch_0_Thresholding_Batcc5D_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccIz.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccIz_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccIz_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccIz(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccIz_rom Thresholding_Batch_0_Thresholding_BatccIz_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingDataWidthConverter_Batch_4_0/synth/finn_design_StreamingDataWidthConverter_Batch_4_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingDataWidthConverter_Batch_4:1.0
// IP Revision: 2101301321

(* X_CORE_INFO = "StreamingDataWidthConverter_Batch_4_StreamingDataWidthConverter_Batch_4,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingDataWidthConverter_Batch_4_0,StreamingDataWidthConverter_Batch_4_StreamingDataWidthConverter_Batch_4,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingDataWidthConverter_Batch_4_0,StreamingDataWidthConverter_Batch_4_StreamingDataWidthConverter_Batch_4,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingDataWidthConverter_Batch_4,x_ipVersion=1.0,x_ipCoreRevision=2101301321,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingDataWidthConverter_Batch_4_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 4, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [31 : 0] out_V_V_TDATA;

  StreamingDataWidthConverter_Batch_4_StreamingDataWidthConverter_Batch_4 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_1_wstrm_0/synth/finn_design_StreamingFCLayer_Batch_1_wstrm_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:user:memstream:1.0
// IP Revision: 5

(* X_CORE_INFO = "memstream,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_1_wstrm_0,memstream,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_1_wstrm_0,memstream,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=user,x_ipName=memstream,x_ipVersion=1.0,x_ipCoreRevision=5,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED,CONFIG_EN=true,NSTREAMS=1,MEM_DEPTH=36864,MEM_WIDTH=64,MEM_INIT=/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/,RAM_STYLE=auto,STRM0_WIDTH=64,STRM1_WIDTH=32,STRM2_WIDTH=32,STRM3_WIDTH=32,STRM4_WIDTH=32,STRM5_WIDTH=32,STR\
M0_DEPTH=36864,STRM1_DEPTH=2304,STRM2_DEPTH=2304,STRM3_DEPTH=2304,STRM4_DEPTH=2304,STRM5_DEPTH=2304,STRM0_OFFSET=0,STRM1_OFFSET=2304,STRM2_OFFSET=4608,STRM3_OFFSET=6912,STRM4_OFFSET=9216,STRM5_OFFSET=11520,AXILITE_ADDR_WIDTH=19}" *)
(* IP_DEFINITION_SOURCE = "package_project" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_1_wstrm_0 (
  aclk,
  aresetn,
  awready,
  awvalid,
  awaddr,
  awprot,
  wready,
  wvalid,
  wdata,
  wstrb,
  bready,
  bvalid,
  bresp,
  arready,
  arvalid,
  araddr,
  arprot,
  rready,
  rvalid,
  rresp,
  rdata,
  m_axis_0_tready,
  m_axis_0_tvalid,
  m_axis_0_tdata
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aclk, ASSOCIATED_BUSIF m_axis_0:m_axis_1:m_axis_2:m_axis_3:m_axis_4:m_axis_5:s_axilite, ASSOCIATED_RESET aresetn, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 aclk CLK" *)
input wire aclk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aresetn, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 aresetn RST" *)
input wire aresetn;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWREADY" *)
output wire awready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWVALID" *)
input wire awvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWADDR" *)
input wire [18 : 0] awaddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWPROT" *)
input wire [2 : 0] awprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WREADY" *)
output wire wready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WVALID" *)
input wire wvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WDATA" *)
input wire [31 : 0] wdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WSTRB" *)
input wire [3 : 0] wstrb;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BREADY" *)
input wire bready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BVALID" *)
output wire bvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BRESP" *)
output wire [1 : 0] bresp;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARREADY" *)
output wire arready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARVALID" *)
input wire arvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARADDR" *)
input wire [18 : 0] araddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARPROT" *)
input wire [2 : 0] arprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RREADY" *)
input wire rready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RVALID" *)
output wire rvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RRESP" *)
output wire [1 : 0] rresp;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axilite, DATA_WIDTH 32, PROTOCOL AXI4LITE, FREQ_HZ 100000000.000000, ID_WIDTH 0, ADDR_WIDTH 19, AWUSER_WIDTH 0, ARUSER_WIDTH 0, WUSER_WIDTH 0, RUSER_WIDTH 0, BUSER_WIDTH 0, READ_WRITE_MODE READ_WRITE, HAS_BURST 0, HAS_LOCK 0, HAS_PROT 1, HAS_CACHE 0, HAS_QOS 0, HAS_REGION 0, HAS_WSTRB 1, HAS_BRESP 1, HAS_RRESP 1, SUPPORTS_NARROW_BURST 0, NUM_READ_OUTSTANDING 1, NUM_WRITE_OUTSTANDING 1, MAX_BURST_LENGTH 1, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, NUM_READ_THREADS 1, NUM_W\
RITE_THREADS 1, RUSER_BITS_PER_BYTE 0, WUSER_BITS_PER_BYTE 0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RDATA" *)
output wire [31 : 0] rdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TREADY" *)
input wire m_axis_0_tready;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TVALID" *)
output wire m_axis_0_tvalid;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME m_axis_0, TDATA_NUM_BYTES 8, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TDATA" *)
output wire [63 : 0] m_axis_0_tdata;

  memstream #(
    .CONFIG_EN(1'B1),
    .NSTREAMS(1),
    .MEM_DEPTH(36864),
    .MEM_WIDTH(64),
    .MEM_INIT("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/"),
    .RAM_STYLE("auto"),
    .STRM0_WIDTH(64),
    .STRM1_WIDTH(32),
    .STRM2_WIDTH(32),
    .STRM3_WIDTH(32),
    .STRM4_WIDTH(32),
    .STRM5_WIDTH(32),
    .STRM0_DEPTH(36864),
    .STRM1_DEPTH(2304),
    .STRM2_DEPTH(2304),
    .STRM3_DEPTH(2304),
    .STRM4_DEPTH(2304),
    .STRM5_DEPTH(2304),
    .STRM0_OFFSET(0),
    .STRM1_OFFSET(2304),
    .STRM2_OFFSET(4608),
    .STRM3_OFFSET(6912),
    .STRM4_OFFSET(9216),
    .STRM5_OFFSET(11520),
    .AXILITE_ADDR_WIDTH(19)
  ) inst (
    .aclk(aclk),
    .aresetn(aresetn),
    .awready(awready),
    .awvalid(awvalid),
    .awaddr(awaddr),
    .awprot(awprot),
    .wready(wready),
    .wvalid(wvalid),
    .wdata(wdata),
    .wstrb(wstrb),
    .bready(bready),
    .bvalid(bvalid),
    .bresp(bresp),
    .arready(arready),
    .arvalid(arvalid),
    .araddr(araddr),
    .arprot(arprot),
    .rready(rready),
    .rvalid(rvalid),
    .rresp(rresp),
    .rdata(rdata),
    .m_axis_0_afull(1'B0),
    .m_axis_0_tready(m_axis_0_tready),
    .m_axis_0_tvalid(m_axis_0_tvalid),
    .m_axis_0_tdata(m_axis_0_tdata),
    .m_axis_1_afull(1'B0),
    .m_axis_1_tready(1'B1),
    .m_axis_1_tvalid(),
    .m_axis_1_tdata(),
    .m_axis_2_afull(1'B0),
    .m_axis_2_tready(1'B1),
    .m_axis_2_tvalid(),
    .m_axis_2_tdata(),
    .m_axis_3_afull(1'B0),
    .m_axis_3_tready(1'B1),
    .m_axis_3_tvalid(),
    .m_axis_3_tdata(),
    .m_axis_4_afull(1'B0),
    .m_axis_4_tready(1'B1),
    .m_axis_4_tvalid(),
    .m_axis_4_tdata(),
    .m_axis_5_afull(1'B0),
    .m_axis_5_tready(1'B1),
    .m_axis_5_tvalid(),
    .m_axis_5_tdata()
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActrcU.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActrcU_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActrcU_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActrcU(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActrcU_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActrcU_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_StreamingFCLayer_Batch_2.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingFCLayer_Batch_2_StreamingFCLayer_Batch_2,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.115000,HLS_SYN_LAT=129607,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=1564,HLS_SYN_LUT=3556,HLS_VERSION=2020_1_1}" *)

module StreamingFCLayer_Batch_2_StreamingFCLayer_Batch_2 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        weights_V_V_TDATA,
        weights_V_V_TVALID,
        weights_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [23:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
input  [47:0] weights_V_V_TDATA;
input   weights_V_V_TVALID;
output   weights_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;
reg weights_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_Matrix_Vector_Activa_fu_140_ap_start;
wire    grp_Matrix_Vector_Activa_fu_140_ap_done;
wire    grp_Matrix_Vector_Activa_fu_140_ap_idle;
wire    grp_Matrix_Vector_Activa_fu_140_ap_ready;
wire    grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY;
wire   [15:0] grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA;
wire    grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID;
wire    grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY;
wire    grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY;
reg    grp_Matrix_Vector_Activa_fu_140_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [23:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    regslice_both_weights_V_V_U_apdone_blk;
wire   [47:0] weights_V_V_TDATA_int;
wire    weights_V_V_TVALID_int;
reg    weights_V_V_TREADY_int;
wire    regslice_both_weights_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_Matrix_Vector_Activa_fu_140_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingFCLayer_Batch_2_Matrix_Vector_Activa grp_Matrix_Vector_Activa_fu_140(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_Matrix_Vector_Activa_fu_140_ap_start),
    .ap_done(grp_Matrix_Vector_Activa_fu_140_ap_done),
    .ap_idle(grp_Matrix_Vector_Activa_fu_140_ap_idle),
    .ap_ready(grp_Matrix_Vector_Activa_fu_140_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY),
    .out_V_V_TDATA(grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA),
    .out_V_V_TVALID(grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID),
    .out_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY),
    .weight_V_V_TDATA(weights_V_V_TDATA_int),
    .weight_V_V_TVALID(weights_V_V_TVALID_int),
    .weight_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 24 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 48 ))
regslice_both_weights_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(weights_V_V_TDATA),
    .vld_in(weights_V_V_TVALID),
    .ack_in(regslice_both_weights_V_V_U_ack_in),
    .data_out(weights_V_V_TDATA_int),
    .vld_out(weights_V_V_TVALID_int),
    .ack_out(weights_V_V_TREADY_int),
    .apdone_blk(regslice_both_weights_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA),
    .vld_in(grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b1;
        end else if ((grp_Matrix_Vector_Activa_fu_140_ap_ready == 1'b1)) begin
            grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    if (((regslice_both_weights_V_V_U_ack_in == 1'b1) & (weights_V_V_TVALID == 1'b1))) begin
        weights_V_V_TREADY = 1'b1;
    end else begin
        weights_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        weights_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY;
    end else begin
        weights_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_Matrix_Vector_Activa_fu_140_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_Matrix_Vector_Activa_fu_140_ap_start = grp_Matrix_Vector_Activa_fu_140_ap_start_reg;

assign grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingFCLayer_Batch_2_StreamingFCLayer_Batch_2
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActRg6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActRg6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActRg6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActRg6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActRg6_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActRg6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_4_0/synth/finn_design_StreamingFCLayer_Batch_4_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFCLayer_Batch_4:1.0
// IP Revision: 2101301316

(* X_CORE_INFO = "StreamingFCLayer_Batch_4_StreamingFCLayer_Batch_4,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_4_0,StreamingFCLayer_Batch_4_StreamingFCLayer_Batch_4,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_4_0,StreamingFCLayer_Batch_4_StreamingFCLayer_Batch_4,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFCLayer_Batch_4,x_ipVersion=1.0,x_ipCoreRevision=2101301316,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_4_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  weights_V_V_TVALID,
  weights_V_V_TREADY,
  weights_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:weights_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 4, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [31 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TVALID" *)
input wire weights_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TREADY" *)
output wire weights_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME weights_V_V, TDATA_NUM_BYTES 16, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TDATA" *)
input wire [127 : 0] weights_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;

  StreamingFCLayer_Batch_4_StreamingFCLayer_Batch_4 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .weights_V_V_TVALID(weights_V_V_TVALID),
    .weights_V_V_TREADY(weights_V_V_TREADY),
    .weights_V_V_TDATA(weights_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccnw.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccnw_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccnw_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccnw(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccnw_rom Thresholding_Batch_0_Thresholding_Batccnw_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActKfY.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActKfY_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActKfY_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActKfY(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActKfY_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActKfY_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActlbW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActlbW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActlbW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActlbW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActlbW_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActlbW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcceu.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcceu_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcceu_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcceu(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcceu_rom Thresholding_Batch_0_Thresholding_Batcceu_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actudo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actudo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actudo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actudo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actudo_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actudo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actsc4.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actsc4_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actsc4_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actsc4(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actsc4_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actsc4_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActpcA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActpcA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActpcA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActpcA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActpcA_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActpcA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcncg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_Batcncg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcncg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_Batcncg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_Batcncg_rom Thresholding_Batch_1_Thresholding_Batcncg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcVhK.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcVhK_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcVhK_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcVhK(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcVhK_rom Thresholding_Batch_0_Thresholding_BatcVhK_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActQgW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActQgW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActQgW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActQgW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActQgW_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActQgW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActWhU.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActWhU_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActWhU_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActWhU(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActWhU_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActWhU_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/5192/StreamingFIFO_7.v


module StreamingFIFO_7(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [23:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [23:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(24)
)
StreamingFIFO_7_StreamingFIFO_7
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActGfk.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActGfk_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActGfk_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActGfk(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActGfk_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActGfk_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_3_0/synth/finn_design_StreamingFCLayer_Batch_3_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFCLayer_Batch_2:1.0
// IP Revision: 2101301318

(* X_CORE_INFO = "StreamingFCLayer_Batch_2_StreamingFCLayer_Batch_2,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_3_0,StreamingFCLayer_Batch_2_StreamingFCLayer_Batch_2,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_3_0,StreamingFCLayer_Batch_2_StreamingFCLayer_Batch_2,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFCLayer_Batch_2,x_ipVersion=1.0,x_ipCoreRevision=2101301318,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_3_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  weights_V_V_TVALID,
  weights_V_V_TREADY,
  weights_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:weights_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 3, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [23 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TVALID" *)
input wire weights_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TREADY" *)
output wire weights_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME weights_V_V, TDATA_NUM_BYTES 6, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TDATA" *)
input wire [47 : 0] weights_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;

  StreamingFCLayer_Batch_2_StreamingFCLayer_Batch_2 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .weights_V_V_TVALID(weights_V_V_TVALID),
    .weights_V_V_TREADY(weights_V_V_TREADY),
    .weights_V_V_TDATA(weights_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/209a/hdl/ramb18_wf_dualport.v

/*
 Copyright (c) 2020, Xilinx
 All rights reserved.

 Redistribution and use in source and binary forms, with or without
 modification, are permitted provided that the following conditions are met:

 * Redistributions of source code must retain the above copyright notice, this
   list of conditions and the following disclaimer.

 * Redistributions in binary form must reproduce the above copyright notice,
   this list of conditions and the following disclaimer in the documentation
   and/or other materials provided with the distribution.

 * Neither the name of FINN nor the names of its
   contributors may be used to endorse or promote products derived from
   this software without specific prior written permission.

 THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
 FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
 SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
 CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
 OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

module ramb18_wf_dualport
#(
    parameter ID = 0,
    parameter DWIDTH = 18,
    parameter AWIDTH = 10,
    parameter DEPTH = 2**AWIDTH,
    parameter MEM_INIT = "",
    parameter RAM_STYLE = "auto"
)
(
	input clk,

	input wea,
    input ena,
    input enqa,
	input [AWIDTH-1:0] addra,
	input [DWIDTH-1:0] wdataa,
	output reg [DWIDTH-1:0] rdqa,

	input web,
    input enb,
    input enqb,
	input [AWIDTH-1:0] addrb,
	input [DWIDTH-1:0] wdatab,
	output reg [DWIDTH-1:0] rdqb
);

(* ram_style = RAM_STYLE *) reg [DWIDTH-1:0] mem[0:DEPTH-1];
reg [DWIDTH-1:0] rdataa;
reg [DWIDTH-1:0] rdatab;

`ifdef SYNTHESIS
reg [7:0] idx = ID;
`else
reg [15:0] idx;
`endif

//initialize memory
initial begin
  //note the hacky way of adding a filename memblock_ID.dat to the path provided in MEM_INIT
  //ID can go up to 99
  if (ID < 0 && ID > 99) begin
    $display("ID out of range [0-99]");
    $finish();
  end
	//MEM_INIT path must be terminated by /
  `ifdef SYNTHESIS
  if (ID < 10)
    $readmemh({MEM_INIT,"memblock_",idx+8'd48,".dat"}, mem, 0, DEPTH-1);
  else
    $readmemh({MEM_INIT,"memblock_",(idx/10)+8'd48,(idx%10)+8'd48,".dat"}, mem, 0, DEPTH-1);
  `else
  $sformat(idx,"%0d",ID);
  if (ID < 10)
    $readmemh({MEM_INIT,"memblock_",idx[7:0],".dat"}, mem, 0, DEPTH-1);
  else
    $readmemh({MEM_INIT,"memblock_",idx,".dat"}, mem, 0, DEPTH-1);
  `endif
end

//memory ports, with output pipeline register
always @(posedge clk) begin
    if(ena) begin
        if(wea)
            mem[addra] <= wdataa;
        rdataa <= mem[addra];
    end
    if(enqa)
        rdqa <= rdataa;
end
always @(posedge clk) begin
    if(enb) begin
        if(web)
            mem[addrb] <= wdatab;
        rdatab <= mem[addrb];
    end
    if(enqb)
        rdqb <= rdatab;
end

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActxdS.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActxdS_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActxdS_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActxdS(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActxdS_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActxdS_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActwdI.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActwdI_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActwdI_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActwdI(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActwdI_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActwdI_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActKfY.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActKfY_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActKfY_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActKfY(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActKfY_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActKfY_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc4D.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcc4D_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc4D_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcc4D(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcc4D_rom Thresholding_Batch_0_Thresholding_Batcc4D_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/af90/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdgE.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcdgE_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdgE_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcdgE(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcdgE_rom Thresholding_Batch_0_Thresholding_BatcdgE_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccqw.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccqw_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccqw_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccqw(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccqw_rom Thresholding_Batch_0_Thresholding_Batccqw_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbqm.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbqm_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbqm_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbqm(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbqm_rom Thresholding_Batch_0_Thresholding_Batcbqm_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActpcA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActpcA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActpcA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActpcA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActpcA_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActpcA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/89c3/StreamingFIFO_15.v


module StreamingFIFO_15(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [31:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(32)
)
StreamingFIFO_15_StreamingFIFO_15
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActkbM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActkbM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActkbM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActkbM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActkbM_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActkbM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actudo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actudo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actudo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actudo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actudo_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actudo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbBo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcbBo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbBo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcbBo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcbBo_rom Thresholding_Batch_0_Thresholding_BatcbBo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActEe0.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActEe0_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActEe0_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActEe0(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActEe0_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActEe0_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActOgC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActOgC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActOgC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActOgC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActOgC_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActOgC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/af90/StreamingFIFO_2.v


module StreamingFIFO_2(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(16)
)
StreamingFIFO_2_StreamingFIFO_2
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcmb6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_Batcmb6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcmb6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_Batcmb6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_Batcmb6_rom Thresholding_Batch_1_Thresholding_Batcmb6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_StreamingFCLayer_5jm.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module StreamingFCLayer_Batch_3_StreamingFCLayer_5jm #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH       = 32,
    din5_WIDTH       = 32,
    din6_WIDTH       = 32,
    din7_WIDTH       = 32,
    din8_WIDTH       = 32,
    din9_WIDTH       = 32,
    din10_WIDTH       = 32,
    din11_WIDTH       = 32,
    din12_WIDTH       = 32,
    din13_WIDTH       = 32,
    din14_WIDTH       = 32,
    din15_WIDTH       = 32,
    din16_WIDTH       = 32,
    din17_WIDTH       = 32,
    din18_WIDTH       = 32,
    din19_WIDTH       = 32,
    din20_WIDTH       = 32,
    din21_WIDTH       = 32,
    din22_WIDTH       = 32,
    din23_WIDTH       = 32,
    din24_WIDTH       = 32,
    din25_WIDTH       = 32,
    din26_WIDTH       = 32,
    din27_WIDTH       = 32,
    din28_WIDTH       = 32,
    din29_WIDTH       = 32,
    din30_WIDTH       = 32,
    din31_WIDTH       = 32,
    din32_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [31 : 0]     din0,
    input  [31 : 0]     din1,
    input  [31 : 0]     din2,
    input  [31 : 0]     din3,
    input  [31 : 0]     din4,
    input  [31 : 0]     din5,
    input  [31 : 0]     din6,
    input  [31 : 0]     din7,
    input  [31 : 0]     din8,
    input  [31 : 0]     din9,
    input  [31 : 0]     din10,
    input  [31 : 0]     din11,
    input  [31 : 0]     din12,
    input  [31 : 0]     din13,
    input  [31 : 0]     din14,
    input  [31 : 0]     din15,
    input  [31 : 0]     din16,
    input  [31 : 0]     din17,
    input  [31 : 0]     din18,
    input  [31 : 0]     din19,
    input  [31 : 0]     din20,
    input  [31 : 0]     din21,
    input  [31 : 0]     din22,
    input  [31 : 0]     din23,
    input  [31 : 0]     din24,
    input  [31 : 0]     din25,
    input  [31 : 0]     din26,
    input  [31 : 0]     din27,
    input  [31 : 0]     din28,
    input  [31 : 0]     din29,
    input  [31 : 0]     din30,
    input  [31 : 0]     din31,
    input  [4 : 0]    din32,
    output [31 : 0]   dout);

// puts internal signals
wire [4 : 0]     sel;
// level 1 signals
wire [31 : 0]         mux_1_0;
wire [31 : 0]         mux_1_1;
wire [31 : 0]         mux_1_2;
wire [31 : 0]         mux_1_3;
wire [31 : 0]         mux_1_4;
wire [31 : 0]         mux_1_5;
wire [31 : 0]         mux_1_6;
wire [31 : 0]         mux_1_7;
wire [31 : 0]         mux_1_8;
wire [31 : 0]         mux_1_9;
wire [31 : 0]         mux_1_10;
wire [31 : 0]         mux_1_11;
wire [31 : 0]         mux_1_12;
wire [31 : 0]         mux_1_13;
wire [31 : 0]         mux_1_14;
wire [31 : 0]         mux_1_15;
// level 2 signals
wire [31 : 0]         mux_2_0;
wire [31 : 0]         mux_2_1;
wire [31 : 0]         mux_2_2;
wire [31 : 0]         mux_2_3;
wire [31 : 0]         mux_2_4;
wire [31 : 0]         mux_2_5;
wire [31 : 0]         mux_2_6;
wire [31 : 0]         mux_2_7;
// level 3 signals
wire [31 : 0]         mux_3_0;
wire [31 : 0]         mux_3_1;
wire [31 : 0]         mux_3_2;
wire [31 : 0]         mux_3_3;
// level 4 signals
wire [31 : 0]         mux_4_0;
wire [31 : 0]         mux_4_1;
// level 5 signals
wire [31 : 0]         mux_5_0;

assign sel = din32;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;
assign mux_1_2 = (sel[0] == 0)? din4 : din5;
assign mux_1_3 = (sel[0] == 0)? din6 : din7;
assign mux_1_4 = (sel[0] == 0)? din8 : din9;
assign mux_1_5 = (sel[0] == 0)? din10 : din11;
assign mux_1_6 = (sel[0] == 0)? din12 : din13;
assign mux_1_7 = (sel[0] == 0)? din14 : din15;
assign mux_1_8 = (sel[0] == 0)? din16 : din17;
assign mux_1_9 = (sel[0] == 0)? din18 : din19;
assign mux_1_10 = (sel[0] == 0)? din20 : din21;
assign mux_1_11 = (sel[0] == 0)? din22 : din23;
assign mux_1_12 = (sel[0] == 0)? din24 : din25;
assign mux_1_13 = (sel[0] == 0)? din26 : din27;
assign mux_1_14 = (sel[0] == 0)? din28 : din29;
assign mux_1_15 = (sel[0] == 0)? din30 : din31;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;
assign mux_2_1 = (sel[1] == 0)? mux_1_2 : mux_1_3;
assign mux_2_2 = (sel[1] == 0)? mux_1_4 : mux_1_5;
assign mux_2_3 = (sel[1] == 0)? mux_1_6 : mux_1_7;
assign mux_2_4 = (sel[1] == 0)? mux_1_8 : mux_1_9;
assign mux_2_5 = (sel[1] == 0)? mux_1_10 : mux_1_11;
assign mux_2_6 = (sel[1] == 0)? mux_1_12 : mux_1_13;
assign mux_2_7 = (sel[1] == 0)? mux_1_14 : mux_1_15;

// Generate level 3 logic
assign mux_3_0 = (sel[2] == 0)? mux_2_0 : mux_2_1;
assign mux_3_1 = (sel[2] == 0)? mux_2_2 : mux_2_3;
assign mux_3_2 = (sel[2] == 0)? mux_2_4 : mux_2_5;
assign mux_3_3 = (sel[2] == 0)? mux_2_6 : mux_2_7;

// Generate level 4 logic
assign mux_4_0 = (sel[3] == 0)? mux_3_0 : mux_3_1;
assign mux_4_1 = (sel[3] == 0)? mux_3_2 : mux_3_3;

// Generate level 5 logic
assign mux_5_0 = (sel[4] == 0)? mux_4_0 : mux_4_1;

// output logic
assign dout = mux_5_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActeOg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActeOg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActeOg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActeOg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActeOg_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActeOg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_10_0/synth/finn_design_StreamingFIFO_10_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_10:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_10,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_10_0,StreamingFIFO_10,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_10_0,StreamingFIFO_10,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_10,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_10_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_10 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/bc91/hdl/verilog/StreamingFCLayer_Batch_6_StreamingFCLayer_cud.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

(* use_dsp = "no" *) module StreamingFCLayer_Batch_6_StreamingFCLayer_cud_Mul_LUT_0(a, b, p);
input[4 - 1 : 0] a; 
input[4 - 1 : 0] b; 
output[8 - 1 : 0] p;

assign p = $signed(a) * $signed(b);
endmodule
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_6_StreamingFCLayer_cud(
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



StreamingFCLayer_Batch_6_StreamingFCLayer_cud_Mul_LUT_0 StreamingFCLayer_Batch_6_StreamingFCLayer_cud_Mul_LUT_0_U(
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcudo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcudo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 5;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcudo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcudo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd5;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcudo_rom Thresholding_Batch_0_Thresholding_Batcudo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actvdy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actvdy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actvdy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actvdy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actvdy_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actvdy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actg8j.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actg8j_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actg8j_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actg8j(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actg8j_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actg8j_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/f5c4/StreamingFIFO_11.v


module StreamingFIFO_11(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(16)
)
StreamingFIFO_11_StreamingFIFO_11
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccQA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccQA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccQA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccQA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccQA_rom Thresholding_Batch_0_Thresholding_BatccQA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActThq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActThq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActThq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActThq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActThq_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActThq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbml.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbml_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbml_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbml(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbml_rom Thresholding_Batch_0_Thresholding_Batcbml_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActUhA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActUhA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActUhA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActUhA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActUhA_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActUhA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8799/StreamingFIFO_16.v


module StreamingFIFO_16(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [7:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(8)
)
StreamingFIFO_16_StreamingFIFO_16
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actocq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actocq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actocq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actocq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actocq_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actocq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Act1iI.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Act1iI_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Act1iI_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Act1iI(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Act1iI_rom StreamingFCLayer_Batch_4_Matrix_Vector_Act1iI_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActeOg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActeOg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActeOg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActeOg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActeOg_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActeOg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActShg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActShg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActShg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActShg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActShg_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActShg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActBew.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActBew_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActBew_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActBew(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActBew_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActBew_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccux.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccux_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccux_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccux(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccux_rom Thresholding_Batch_0_Thresholding_Batccux_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/209a/hdl/memstream_multiblock.v

/*
 Copyright (c) 2020, Xilinx
 All rights reserved.

 Redistribution and use in source and binary forms, with or without
 modification, are permitted provided that the following conditions are met:

 * Redistributions of source code must retain the above copyright notice, this
   list of conditions and the following disclaimer.

 * Redistributions in binary form must reproduce the above copyright notice,
   this list of conditions and the following disclaimer in the documentation
   and/or other materials provided with the distribution.

 * Neither the name of FINN nor the names of its
   contributors may be used to endorse or promote products derived from
   this software without specific prior written permission.

 THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
 FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
 SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
 CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
 OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

module memstream_multiblock
#(
//parameters to enable/disable axi-mm, set number of streams, set readmemh for memory, set per-stream offsets in memory, set per-stream widths
    parameter CONFIG_EN = 1,
    parameter NSTREAMS = 6,//1 up to 6

    parameter MEM_DEPTH = 13824,
    parameter MEM_WIDTH = 32,
    parameter MEM_INIT = "./",
    parameter RAM_STYLE = "auto",

    //widths per stream
	parameter STRM0_WIDTH = 32,
	parameter STRM1_WIDTH = 32,
	parameter STRM2_WIDTH = 32,
	parameter STRM3_WIDTH = 32,
	parameter STRM4_WIDTH = 32,
	parameter STRM5_WIDTH = 32,

	//depths per stream
	parameter STRM0_DEPTH = 2304,
	parameter STRM1_DEPTH = 2304,
	parameter STRM2_DEPTH = 2304,
	parameter STRM3_DEPTH = 2304,
	parameter STRM4_DEPTH = 2304,
	parameter STRM5_DEPTH = 2304,

	//offsets for each stream
	parameter STRM0_OFFSET = 0,
	parameter STRM1_OFFSET = 2304,
	parameter STRM2_OFFSET = 4608,
	parameter STRM3_OFFSET = 6912,
	parameter STRM4_OFFSET = 9216,
	parameter STRM5_OFFSET = 11520
)

(
    input aclk,
    input aresetn,

    //optional configuration interface compatible with ap_memory
	input [31:0] config_address,
	input config_ce,
	input config_we,
	input [31:0] config_d0,
	output [31:0] config_q0,
    output config_rack,

    //multiple output AXI Streams, TDATA width rounded to multiple of 8 bits
    input m_axis_0_afull,
    input m_axis_0_tready,
    output m_axis_0_tvalid,
    output [((STRM0_WIDTH+7)/8)*8-1:0] m_axis_0_tdata,

    input m_axis_1_afull,
    input m_axis_1_tready,
    output m_axis_1_tvalid,
    output [((STRM1_WIDTH+7)/8)*8-1:0] m_axis_1_tdata,

    input m_axis_2_afull,
    input m_axis_2_tready,
    output m_axis_2_tvalid,
    output [((STRM2_WIDTH+7)/8)*8-1:0] m_axis_2_tdata,

    input m_axis_3_afull,
    input m_axis_3_tready,
    output m_axis_3_tvalid,
    output [((STRM3_WIDTH+7)/8)*8-1:0] m_axis_3_tdata,

    input m_axis_4_afull,
    input m_axis_4_tready,
    output m_axis_4_tvalid,
    output [((STRM4_WIDTH+7)/8)*8-1:0] m_axis_4_tdata,

    input m_axis_5_afull,
    input m_axis_5_tready,
    output m_axis_5_tvalid,
    output [((STRM5_WIDTH+7)/8)*8-1:0] m_axis_5_tdata


);

//calculate number of RAMB18 blocks we need depth-wise
localparam NMEMBLOCKS = (MEM_DEPTH+1023) / 1024; //ceil(MEM_DEPTH/1024)

//calculate width of address for each block
localparam BLOCKADRWIDTH = NMEMBLOCKS > 1 ? 10 : $clog2(MEM_DEPTH);

//determine whether a stream needs to multiplex between memory blocks
localparam STRM0_MUX = ((STRM0_OFFSET/1024) != ((STRM0_OFFSET+STRM0_DEPTH)/1024));
localparam STRM1_MUX = ((STRM1_OFFSET/1024) != ((STRM1_OFFSET+STRM1_DEPTH)/1024));
localparam STRM2_MUX = ((STRM2_OFFSET/1024) != ((STRM2_OFFSET+STRM2_DEPTH)/1024));
localparam STRM3_MUX = ((STRM3_OFFSET/1024) != ((STRM3_OFFSET+STRM3_DEPTH)/1024));
localparam STRM4_MUX = ((STRM4_OFFSET/1024) != ((STRM4_OFFSET+STRM4_DEPTH)/1024));
localparam STRM5_MUX = ((STRM5_OFFSET/1024) != ((STRM5_OFFSET+STRM5_DEPTH)/1024));

//determine what the base block of each stream is
localparam STRM0_BLOCK = (STRM0_OFFSET/1024);
localparam STRM1_BLOCK = (STRM1_OFFSET/1024);
localparam STRM2_BLOCK = (STRM2_OFFSET/1024);
localparam STRM3_BLOCK = (STRM3_OFFSET/1024);
localparam STRM4_BLOCK = (STRM4_OFFSET/1024);
localparam STRM5_BLOCK = (STRM5_OFFSET/1024);

//determine what the end block of each stream is
localparam STRM0_END_BLOCK = ((STRM0_OFFSET+STRM0_DEPTH-1)/1024);
localparam STRM1_END_BLOCK = ((STRM1_OFFSET+STRM1_DEPTH-1)/1024);
localparam STRM2_END_BLOCK = ((STRM2_OFFSET+STRM2_DEPTH-1)/1024);
localparam STRM3_END_BLOCK = ((STRM3_OFFSET+STRM3_DEPTH-1)/1024);
localparam STRM4_END_BLOCK = ((STRM4_OFFSET+STRM4_DEPTH-1)/1024);
localparam STRM5_END_BLOCK = ((STRM5_OFFSET+STRM5_DEPTH-1)/1024);

//determine the number of blocks spanned by each stream
localparam STRM0_NBLOCKS = STRM0_END_BLOCK - STRM0_BLOCK + 1;
localparam STRM1_NBLOCKS = STRM1_END_BLOCK - STRM1_BLOCK + 1;
localparam STRM2_NBLOCKS = STRM2_END_BLOCK - STRM2_BLOCK + 1;
localparam STRM3_NBLOCKS = STRM3_END_BLOCK - STRM3_BLOCK + 1;
localparam STRM4_NBLOCKS = STRM4_END_BLOCK - STRM4_BLOCK + 1;
localparam STRM5_NBLOCKS = STRM5_END_BLOCK - STRM5_BLOCK + 1;

//TODO: check that memory width is equal to the widest stream
//TODO: check that the stream depths and offsets make sense, and that the memory depth is sufficient (or calculate depth here?)
initial begin
    if((NSTREAMS < 1) | (NSTREAMS > 6)) begin
        $display("Invalid setting for NSTREAMS, please set in range [1,6]");
        $finish();
    end
end

//invert reset
wire rst;
assign rst = ~aresetn;

//WARNING: pipeline depth is larger than the number of streams per port so we have in-flight writes that may see not-ready when they get executed
//solution: use prog-full to make sure we have an equal number of free slots in the stream to the read pipeline depth

reg [$clog2(MEM_DEPTH)-1:0] strm0_addr = STRM0_OFFSET;
reg [$clog2(MEM_DEPTH)-1:0] strm1_addr = STRM1_OFFSET;
reg [$clog2(MEM_DEPTH)-1:0] strm2_addr = STRM2_OFFSET;
reg [$clog2(MEM_DEPTH)-1:0] strm3_addr = STRM3_OFFSET;
reg [$clog2(MEM_DEPTH)-1:0] strm4_addr = STRM4_OFFSET;
reg [$clog2(MEM_DEPTH)-1:0] strm5_addr = STRM5_OFFSET;

reg strm0_incr_en;
reg strm1_incr_en;
reg strm2_incr_en;
reg strm3_incr_en;
reg strm4_incr_en;
reg strm5_incr_en;

wire strm0_rst;
wire strm1_rst;
wire strm2_rst;
wire strm3_rst;
wire strm4_rst;
wire strm5_rst;

reg strm0_ready;
reg strm1_ready;
reg strm2_ready;
reg strm3_ready;
reg strm4_ready;
reg strm5_ready;

//arbiter: work on one stream at a time
//multiplex each port between (up to) half of the streams
reg [1:0] current_stream_porta = 0;
reg [1:0] current_stream_portb = 0;

always @(posedge aclk) begin
    if(rst)
        current_stream_porta <= 0;
    else case(current_stream_porta)
        0: current_stream_porta <= strm2_ready ? 1 : strm4_ready ? 2 : 0;
        1: current_stream_porta <= strm4_ready ? 2 : strm0_ready ? 0 : 1;
        2: current_stream_porta <= strm0_ready ? 0 : strm2_ready ? 1 : 2;
    endcase
    if(rst)
        current_stream_portb <= 0;
    else case(current_stream_portb)
        0: current_stream_portb <= strm3_ready ? 1 : strm5_ready ? 2 : 0;
        1: current_stream_portb <= strm5_ready ? 2 : strm1_ready ? 0 : 1;
        2: current_stream_portb <= strm1_ready ? 0 : strm3_ready ? 1 : 2;
    endcase
end

always @(posedge aclk) begin
    if(rst) begin
        strm0_incr_en <= 0;
        strm1_incr_en <= 0;
        strm2_incr_en <= 0;
        strm3_incr_en <= 0;
        strm4_incr_en <= 0;
        strm5_incr_en <= 0;
    end else begin
        strm0_incr_en <= (current_stream_porta == 0) & strm0_ready;
        strm1_incr_en <= (current_stream_portb == 0) & strm1_ready;
        strm2_incr_en <= (current_stream_porta == 1) & strm2_ready;
        strm3_incr_en <= (current_stream_portb == 1) & strm3_ready;
        strm4_incr_en <= (current_stream_porta == 2) & strm4_ready;
        strm5_incr_en <= (current_stream_portb == 2) & strm5_ready;
    end
end

assign strm0_rst = strm0_incr_en & (strm0_addr == (STRM0_OFFSET + STRM0_DEPTH-1));
assign strm1_rst = strm1_incr_en & (strm1_addr == (STRM1_OFFSET + STRM1_DEPTH-1));
assign strm2_rst = strm2_incr_en & (strm2_addr == (STRM2_OFFSET + STRM2_DEPTH-1));
assign strm3_rst = strm3_incr_en & (strm3_addr == (STRM3_OFFSET + STRM3_DEPTH-1));
assign strm4_rst = strm4_incr_en & (strm4_addr == (STRM4_OFFSET + STRM4_DEPTH-1));
assign strm5_rst = strm5_incr_en & (strm5_addr == (STRM5_OFFSET + STRM5_DEPTH-1));

always @(posedge aclk) begin
    strm0_ready <= ~m_axis_0_afull;
    strm1_ready <= ~m_axis_1_afull & (NSTREAMS >= 2);
    strm2_ready <= ~m_axis_2_afull & (NSTREAMS >= 3);
    strm3_ready <= ~m_axis_3_afull & (NSTREAMS >= 4);
    strm4_ready <= ~m_axis_4_afull & (NSTREAMS >= 5);
    strm5_ready <= ~m_axis_5_afull & (NSTREAMS >= 6);
end

//one address counter per stream; more LUTs but keeps routing short and local
always @(posedge aclk) begin
    if(strm0_rst | rst)
        strm0_addr <= STRM0_OFFSET;
    else if(strm0_incr_en)
        strm0_addr <= strm0_addr + 1;
    if(strm1_rst | rst)
        strm1_addr <= STRM1_OFFSET;
    else if(strm1_incr_en)
        strm1_addr <= strm1_addr + 1;
    if(strm2_rst | rst)
        strm2_addr <= STRM2_OFFSET;
    else if(strm2_incr_en)
        strm2_addr <= strm2_addr + 1;
    if(strm3_rst | rst)
        strm3_addr <= STRM3_OFFSET;
    else if(strm3_incr_en)
        strm3_addr <= strm3_addr + 1;
    if(strm4_rst | rst)
        strm4_addr <= STRM4_OFFSET;
    else if(strm4_incr_en)
        strm4_addr <= strm4_addr + 1;
    if(strm5_rst | rst)
        strm5_addr <= STRM5_OFFSET;
    else if(strm5_incr_en)
        strm5_addr <= strm5_addr + 1;
end

reg [$clog2(MEM_DEPTH)-1:0] addra;
wire [MEM_WIDTH*NMEMBLOCKS-1:0] rdqa;

reg [$clog2(MEM_DEPTH)-1:0] addrb;
wire [MEM_WIDTH*NMEMBLOCKS-1:0] rdqb;

wire [NMEMBLOCKS-1:0] we;

reg [1:0] addr_select_porta;
reg [1:0] addr_select_portb;

//multiplex addresses of various streams into address ports of memory
always @(posedge aclk) begin
    addr_select_porta <= current_stream_porta;
    case(addr_select_porta)
        0: addra <= strm0_addr;
        1: addra <= strm2_addr;
        2: addra <= strm4_addr;
    endcase
    addr_select_portb <= current_stream_portb;
    case(addr_select_portb)
        0: addrb <= strm1_addr;
        1: addrb <= strm3_addr;
        2: addrb <= strm5_addr;
    endcase
end

genvar g;
generate for(g=0; g<NMEMBLOCKS; g=g+1) begin: blockports

assign we[g] = (CONFIG_EN == 1) & config_ce & config_we & (config_address[31:BLOCKADRWIDTH] == g);

ramb18_wf_dualport
#(
    .ID(g),
	.DWIDTH(MEM_WIDTH),
	.AWIDTH(BLOCKADRWIDTH),
	.MEM_INIT(MEM_INIT),
  .RAM_STYLE(RAM_STYLE)
)
ram
(
	.clk(aclk),

	.wea(we[g]),
    .ena(1'b1),
    .enqa(1'b1),
	.addra(we[g] ? config_address[BLOCKADRWIDTH-1:0] : addra[BLOCKADRWIDTH-1:0]),
	.wdataa(config_d0),
	.rdqa(rdqa[(g+1)*MEM_WIDTH-1:g*MEM_WIDTH]),

	.web(1'b0),
    .enb(1'b1),
    .enqb(1'b1),
	.addrb(addrb[BLOCKADRWIDTH-1:0]),
	.wdatab('d0),
	.rdqb(rdqb[(g+1)*MEM_WIDTH-1:g*MEM_WIDTH])
);

end
endgenerate

integer i;

generate if(NMEMBLOCKS > 1) begin: multiblock

wire [MEM_WIDTH-1:0] rdqmux[5:0];

reg [$clog2(MEM_DEPTH)-BLOCKADRWIDTH-1:0] rdblocka[2:0];
reg [$clog2(MEM_DEPTH)-BLOCKADRWIDTH-1:0] rdblockb[2:0];

always @(posedge aclk) begin
    rdblocka[0] <= addra[$clog2(MEM_DEPTH)-1:BLOCKADRWIDTH];
    rdblockb[0] <= addrb[$clog2(MEM_DEPTH)-1:BLOCKADRWIDTH];
    for(i=0; i<2; i=i+1) begin
		rdblocka[i+1] <= rdblocka[i];
		rdblockb[i+1] <= rdblockb[i];
    end
end

if(NSTREAMS >= 1) begin: en_strm0
	if(STRM0_MUX == 1) begin: mux0
		mux #(STRM0_NBLOCKS, MEM_WIDTH) m(rdqa[(STRM0_BLOCK+STRM0_NBLOCKS)*MEM_WIDTH-1:STRM0_BLOCK*MEM_WIDTH],rdqmux[0],rdblocka[1] - STRM0_BLOCK);
	end else begin: nomux0
		assign rdqmux[0] = rdqa[(STRM0_BLOCK+1)*MEM_WIDTH-1:STRM0_BLOCK*MEM_WIDTH];
	end
	assign m_axis_0_tdata = rdqmux[0][STRM0_WIDTH-1:0];
end

if(NSTREAMS >= 2) begin: en_strm1
	if(STRM1_MUX == 1) begin: mux1
		mux #(STRM1_NBLOCKS, MEM_WIDTH) m(rdqb[(STRM1_BLOCK+STRM1_NBLOCKS)*MEM_WIDTH-1:STRM1_BLOCK*MEM_WIDTH],rdqmux[1],rdblockb[1] - STRM1_BLOCK);
	end else begin: nomux1
		assign rdqmux[1] = rdqb[(STRM1_BLOCK+1)*MEM_WIDTH-1:STRM1_BLOCK*MEM_WIDTH];
	end
	assign m_axis_1_tdata = rdqmux[1][STRM1_WIDTH-1:0];
end

if(NSTREAMS >= 3) begin: en_strm2
	if(STRM2_MUX == 1) begin: mux2
		mux #(STRM2_NBLOCKS, MEM_WIDTH) m(rdqa[(STRM2_BLOCK+STRM2_NBLOCKS)*MEM_WIDTH-1:STRM2_BLOCK*MEM_WIDTH],rdqmux[2],rdblocka[1] - STRM2_BLOCK);
	end else begin: nomux2
		assign rdqmux[2] = rdqa[(STRM2_BLOCK+1)*MEM_WIDTH-1:STRM2_BLOCK*MEM_WIDTH];
	end
	assign m_axis_2_tdata = rdqmux[2][STRM2_WIDTH-1:0];
end

if(NSTREAMS >= 4) begin: en_strm3
	if(STRM3_MUX == 1) begin: mux3
		mux #(STRM3_NBLOCKS, MEM_WIDTH) m(rdqb[(STRM3_BLOCK+STRM3_NBLOCKS)*MEM_WIDTH-1:STRM3_BLOCK*MEM_WIDTH],rdqmux[3],rdblockb[1] - STRM3_BLOCK);
	end else begin: nomux3
		assign rdqmux[3] = rdqb[(STRM3_BLOCK+1)*MEM_WIDTH-1:STRM3_BLOCK*MEM_WIDTH];
	end
	assign m_axis_3_tdata = rdqmux[3][STRM3_WIDTH-1:0];
end

if(NSTREAMS >= 5) begin: en_strm4
	if(STRM4_MUX == 1) begin: mux4
		mux #(STRM4_NBLOCKS, MEM_WIDTH) m(rdqa[(STRM4_BLOCK+STRM4_NBLOCKS)*MEM_WIDTH-1:STRM4_BLOCK*MEM_WIDTH],rdqmux[4],rdblocka[1] - STRM4_BLOCK);
	end else begin: nomux4
		assign rdqmux[4] = rdqa[(STRM4_BLOCK+1)*MEM_WIDTH-1:STRM4_BLOCK*MEM_WIDTH];
	end
	assign m_axis_4_tdata = rdqmux[4][STRM4_WIDTH-1:0];
end

if(NSTREAMS >= 6) begin: en_strm5
	if(STRM5_MUX == 1) begin: mux5
		mux #(STRM5_NBLOCKS, MEM_WIDTH) m(rdqb[(STRM5_BLOCK+STRM5_NBLOCKS)*MEM_WIDTH-1:STRM5_BLOCK*MEM_WIDTH],rdqmux[5],rdblockb[1] - STRM5_BLOCK);
	end else begin: nomux5
		assign rdqmux[5] = rdqb[(STRM5_BLOCK+1)*MEM_WIDTH-1:STRM5_BLOCK*MEM_WIDTH];
	end
	assign m_axis_5_tdata = rdqmux[5][STRM5_WIDTH-1:0];
end

end else begin: singleblock

if(NSTREAMS >= 1) begin: en_strm0_direct
    assign m_axis_0_tdata = rdqa[STRM0_WIDTH-1:0];
end
if(NSTREAMS >= 2) begin: en_strm1_direct
	assign m_axis_1_tdata = rdqb[STRM1_WIDTH-1:0];
end
if(NSTREAMS >= 3) begin: en_strm2_direct
	assign m_axis_2_tdata = rdqa[STRM2_WIDTH-1:0];
end
if(NSTREAMS >= 4) begin: en_strm3_direct
	assign m_axis_3_tdata = rdqb[STRM3_WIDTH-1:0];
end
if(NSTREAMS >= 5) begin: en_strm4_direct
	assign m_axis_4_tdata = rdqa[STRM4_WIDTH-1:0];
end
if(NSTREAMS >= 6) begin: en_strm5_direct
	assign m_axis_5_tdata = rdqb[STRM5_WIDTH-1:0];
end

end
endgenerate

//output to AXI Streams
reg tvalid_pipe0[2:0];
reg tvalid_pipe1[2:0];
reg tvalid_pipe2[2:0];
reg tvalid_pipe3[2:0];
reg tvalid_pipe4[2:0];
reg tvalid_pipe5[2:0];

assign m_axis_0_tvalid = tvalid_pipe0[2];
assign m_axis_1_tvalid = tvalid_pipe1[2];
assign m_axis_2_tvalid = tvalid_pipe2[2];
assign m_axis_3_tvalid = tvalid_pipe3[2];
assign m_axis_4_tvalid = tvalid_pipe4[2];
assign m_axis_5_tvalid = tvalid_pipe5[2];


always @(posedge aclk) begin
    tvalid_pipe0[0] <= strm0_incr_en;
    tvalid_pipe1[0] <= strm1_incr_en;
    tvalid_pipe2[0] <= strm2_incr_en;
    tvalid_pipe3[0] <= strm3_incr_en;
    tvalid_pipe4[0] <= strm4_incr_en;
    tvalid_pipe5[0] <= strm5_incr_en;
    for(i=0; i<2; i=i+1) begin: srl
        tvalid_pipe0[i+1] <= tvalid_pipe0[i];
        tvalid_pipe1[i+1] <= tvalid_pipe1[i];
        tvalid_pipe2[i+1] <= tvalid_pipe2[i];
        tvalid_pipe3[i+1] <= tvalid_pipe3[i];
        tvalid_pipe4[i+1] <= tvalid_pipe4[i];
        tvalid_pipe5[i+1] <= tvalid_pipe5[i];
    end
end

//dummy read, for now
assign config_q0 = 0;
assign config_rack = config_ce & ~config_we;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActdEe.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActdEe_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActdEe_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActdEe(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActdEe_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActdEe_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActCeG.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActCeG_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActCeG_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActCeG(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActCeG_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActCeG_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActMgi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActMgi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActMgi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActMgi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActMgi_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActMgi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcg8j.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_Batcg8j_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcg8j_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_Batcg8j(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_Batcg8j_rom Thresholding_Batch_2_Thresholding_Batcg8j_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_Batchbi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_Batchbi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_Batchbi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_Batchbi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_Batchbi_rom Thresholding_Batch_2_Thresholding_Batchbi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActjbC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActjbC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActjbC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActjbC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActjbC_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActjbC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActdEe.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActdEe_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActdEe_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActdEe(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActdEe_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActdEe_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccKz.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccKz_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccKz_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccKz(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccKz_rom Thresholding_Batch_0_Thresholding_BatccKz_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcJfO.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcJfO_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcJfO_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcJfO(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcJfO_rom Thresholding_Batch_0_Thresholding_BatcJfO_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Act0iy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Act0iy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Act0iy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Act0iy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Act0iy_rom StreamingFCLayer_Batch_2_Matrix_Vector_Act0iy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_18_0/synth/finn_design_StreamingFIFO_18_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_18:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_18,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_18_0,StreamingFIFO_18,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_18_0,StreamingFIFO_18,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_18,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_18_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_18 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActVhK.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActVhK_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActVhK_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActVhK(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActVhK_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActVhK_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActXh4.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActXh4_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActXh4_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActXh4(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActXh4_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActXh4_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccBy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccBy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccBy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccBy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccBy_rom Thresholding_Batch_0_Thresholding_BatccBy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActXh4.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActXh4_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActXh4_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActXh4(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActXh4_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActXh4_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actcud.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actcud_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actcud_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actcud(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actcud_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actcud_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_StreamingFCLayer_Batch_3.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingFCLayer_Batch_3_StreamingFCLayer_Batch_3,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.409000,HLS_SYN_LAT=4104,HLS_SYN_TPT=none,HLS_SYN_MEM=56,HLS_SYN_DSP=0,HLS_SYN_FF=1641,HLS_SYN_LUT=3159,HLS_VERSION=2020_1_1}" *)

module StreamingFCLayer_Batch_3_StreamingFCLayer_Batch_3 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        weights_V_V_TDATA,
        weights_V_V_TVALID,
        weights_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [31:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
input  [127:0] weights_V_V_TDATA;
input   weights_V_V_TVALID;
output   weights_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;
reg weights_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_Matrix_Vector_Activa_fu_140_ap_start;
wire    grp_Matrix_Vector_Activa_fu_140_ap_done;
wire    grp_Matrix_Vector_Activa_fu_140_ap_idle;
wire    grp_Matrix_Vector_Activa_fu_140_ap_ready;
wire    grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY;
wire   [15:0] grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA;
wire    grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID;
wire    grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY;
wire    grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY;
reg    grp_Matrix_Vector_Activa_fu_140_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [31:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    regslice_both_weights_V_V_U_apdone_blk;
wire   [127:0] weights_V_V_TDATA_int;
wire    weights_V_V_TVALID_int;
reg    weights_V_V_TREADY_int;
wire    regslice_both_weights_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_Matrix_Vector_Activa_fu_140_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingFCLayer_Batch_3_Matrix_Vector_Activa grp_Matrix_Vector_Activa_fu_140(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_Matrix_Vector_Activa_fu_140_ap_start),
    .ap_done(grp_Matrix_Vector_Activa_fu_140_ap_done),
    .ap_idle(grp_Matrix_Vector_Activa_fu_140_ap_idle),
    .ap_ready(grp_Matrix_Vector_Activa_fu_140_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY),
    .out_V_V_TDATA(grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA),
    .out_V_V_TVALID(grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID),
    .out_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY),
    .weight_V_V_TDATA(weights_V_V_TDATA_int),
    .weight_V_V_TVALID(weights_V_V_TVALID_int),
    .weight_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 32 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 128 ))
regslice_both_weights_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(weights_V_V_TDATA),
    .vld_in(weights_V_V_TVALID),
    .ack_in(regslice_both_weights_V_V_U_ack_in),
    .data_out(weights_V_V_TDATA_int),
    .vld_out(weights_V_V_TVALID_int),
    .ack_out(weights_V_V_TREADY_int),
    .apdone_blk(regslice_both_weights_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA),
    .vld_in(grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b1;
        end else if ((grp_Matrix_Vector_Activa_fu_140_ap_ready == 1'b1)) begin
            grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    if (((regslice_both_weights_V_V_U_ack_in == 1'b1) & (weights_V_V_TVALID == 1'b1))) begin
        weights_V_V_TREADY = 1'b1;
    end else begin
        weights_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        weights_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY;
    end else begin
        weights_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_Matrix_Vector_Activa_fu_140_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_Matrix_Vector_Activa_fu_140_ap_start = grp_Matrix_Vector_Activa_fu_140_ap_start_reg;

assign grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingFCLayer_Batch_3_StreamingFCLayer_Batch_3
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Acthbi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Acthbi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Acthbi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Acthbi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Acthbi_rom StreamingFCLayer_Batch_2_Matrix_Vector_Acthbi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_LabelSelect_Batch_0_0/synth/finn_design_LabelSelect_Batch_0_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:LabelSelect_Batch_0:1.0
// IP Revision: 2101301315

(* X_CORE_INFO = "LabelSelect_Batch_0_LabelSelect_Batch_0,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_LabelSelect_Batch_0_0,LabelSelect_Batch_0_LabelSelect_Batch_0,{}" *)
(* CORE_GENERATION_INFO = "finn_design_LabelSelect_Batch_0_0,LabelSelect_Batch_0_LabelSelect_Batch_0,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=LabelSelect_Batch_0,x_ipVersion=1.0,x_ipCoreRevision=2101301315,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_LabelSelect_Batch_0_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;

  LabelSelect_Batch_0_LabelSelect_Batch_0 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActJfO.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActJfO_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActJfO_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActJfO(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActJfO_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActJfO_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actncg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actncg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actncg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actncg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actncg_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actncg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActfYi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActfYi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActfYi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActfYi_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActfYi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActNgs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActNgs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActNgs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActNgs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActNgs_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActNgs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actsc4.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actsc4_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actsc4_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actsc4(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actsc4_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actsc4_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/32c2/hdl/verilog/StreamingDataWidthConverter_Batch_5_StreamingDataWidthConverter_Batch_5.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingDataWidthConverter_Batch_5_StreamingDataWidthConverter_Batch_5,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=5.723000,HLS_SYN_LAT=261,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=77,HLS_SYN_LUT=288,HLS_VERSION=2020_1_1}" *)

module StreamingDataWidthConverter_Batch_5_StreamingDataWidthConverter_Batch_5 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_start;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_done;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_idle;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_ready;
wire    grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
wire   [7:0] grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY;
reg    grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [15:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_StreamingDataWidthCo_1_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingDataWidthConverter_Batch_5_StreamingDataWidthCo_1 grp_StreamingDataWidthCo_1_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_StreamingDataWidthCo_1_fu_26_ap_start),
    .ap_done(grp_StreamingDataWidthCo_1_fu_26_ap_done),
    .ap_idle(grp_StreamingDataWidthCo_1_fu_26_ap_idle),
    .ap_ready(grp_StreamingDataWidthCo_1_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .vld_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_StreamingDataWidthCo_1_fu_26_ap_ready == 1'b1)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_StreamingDataWidthCo_1_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_StreamingDataWidthCo_1_fu_26_ap_start = grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;

assign grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingDataWidthConverter_Batch_5_StreamingDataWidthConverter_Batch_5
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actzec.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actzec_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actzec_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actzec(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actzec_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actzec_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccJz.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccJz_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccJz_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccJz(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccJz_rom Thresholding_Batch_0_Thresholding_BatccJz_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actbkb_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actbkb_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actbkb(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actbkb_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actbkb_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActwdI.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActwdI_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActwdI_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActwdI(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActwdI_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActwdI_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/cd9c/hdl/verilog/StreamingFCLayer_Batch_0_StreamingFCLayer_cud.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

(* use_dsp = "no" *) module StreamingFCLayer_Batch_0_StreamingFCLayer_cud_Mul_LUT_0(a, b, p);
input[4 - 1 : 0] a; 
input[4 - 1 : 0] b; 
output[8 - 1 : 0] p;

assign p = $signed(a) * $signed(b);
endmodule
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_0_StreamingFCLayer_cud(
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



StreamingFCLayer_Batch_0_StreamingFCLayer_cud_Mul_LUT_0 StreamingFCLayer_Batch_0_StreamingFCLayer_cud_Mul_LUT_0_U(
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/db73/StreamingFIFO_3.v


module StreamingFIFO_3(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [7:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(8)
)
StreamingFIFO_3_StreamingFIFO_3
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/209a/hdl/memstream.v

/*
 Copyright (c) 2020, Xilinx
 All rights reserved.

 Redistribution and use in source and binary forms, with or without
 modification, are permitted provided that the following conditions are met:

 * Redistributions of source code must retain the above copyright notice, this
   list of conditions and the following disclaimer.

 * Redistributions in binary form must reproduce the above copyright notice,
   this list of conditions and the following disclaimer in the documentation
   and/or other materials provided with the distribution.

 * Neither the name of FINN nor the names of its
   contributors may be used to endorse or promote products derived from
   this software without specific prior written permission.

 THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
 FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
 SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
 CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
 OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

module memstream
#(
//parameters to enable/disable axi-mm, set number of streams, set readmemh for memory, set per-stream offsets in memory, set per-stream widths
    parameter CONFIG_EN = 1,
    parameter NSTREAMS = 6,//1 up to 6

    parameter MEM_DEPTH = 13824,
    parameter MEM_WIDTH = 32,
    parameter MEM_INIT = "./",
    parameter RAM_STYLE = "auto",

    //widths per stream
	parameter STRM0_WIDTH = 32,
	parameter STRM1_WIDTH = 32,
	parameter STRM2_WIDTH = 32,
	parameter STRM3_WIDTH = 32,
	parameter STRM4_WIDTH = 32,
	parameter STRM5_WIDTH = 32,

	//depths per stream
	parameter STRM0_DEPTH = 2304,
	parameter STRM1_DEPTH = 2304,
	parameter STRM2_DEPTH = 2304,
	parameter STRM3_DEPTH = 2304,
	parameter STRM4_DEPTH = 2304,
	parameter STRM5_DEPTH = 2304,

	//offsets for each stream
	parameter STRM0_OFFSET = 0,
	parameter STRM1_OFFSET = 2304,
	parameter STRM2_OFFSET = 4608,
	parameter STRM3_OFFSET = 6912,
	parameter STRM4_OFFSET = 9216,
	parameter STRM5_OFFSET = 11520,

    parameter AXILITE_ADDR_WIDTH = 2+$clog2(MEM_DEPTH*(1<<$clog2((MEM_WIDTH+31)/32)))
)

(
    input aclk,
    input aresetn,

    output awready,
    input                       awvalid,
    input [AXILITE_ADDR_WIDTH-1:0]      awaddr,
    input [2:0]                 awprot,
    //write data
    output                  wready,
    input                       wvalid,
    input [31:0]      wdata,
    input [3:0]  wstrb,
    //burst response
    input                       bready,
    output                  bvalid,
    output [1:0]            bresp,

    //Read channels
    //read address
    output                  arready,
    input                       arvalid,
    input [AXILITE_ADDR_WIDTH-1:0]      araddr,
    input [2:0]                 arprot,
    //read data
    input                       rready,
    output                  rvalid,
    output [1:0]            rresp,
    output [31:0] rdata,

    //multiple output AXI Streams, TDATA width rounded to multiple of 8 bits
    input m_axis_0_afull,
    input m_axis_0_tready,
    output m_axis_0_tvalid,
    output [((STRM0_WIDTH+7)/8)*8-1:0] m_axis_0_tdata,

    input m_axis_1_afull,
    input m_axis_1_tready,
    output m_axis_1_tvalid,
    output [((STRM1_WIDTH+7)/8)*8-1:0] m_axis_1_tdata,

    input m_axis_2_afull,
    input m_axis_2_tready,
    output m_axis_2_tvalid,
    output [((STRM2_WIDTH+7)/8)*8-1:0] m_axis_2_tdata,

    input m_axis_3_afull,
    input m_axis_3_tready,
    output m_axis_3_tvalid,
    output [((STRM3_WIDTH+7)/8)*8-1:0] m_axis_3_tdata,

    input m_axis_4_afull,
    input m_axis_4_tready,
    output m_axis_4_tvalid,
    output [((STRM4_WIDTH+7)/8)*8-1:0] m_axis_4_tdata,

    input m_axis_5_afull,
    input m_axis_5_tready,
    output m_axis_5_tvalid,
    output [((STRM5_WIDTH+7)/8)*8-1:0] m_axis_5_tdata


);

wire [31:0] config_address;
wire config_ce;
wire config_we;
wire config_rack;
wire [MEM_WIDTH-1:0] config_d0;
wire [MEM_WIDTH-1:0] config_q0;

generate
if(NSTREAMS <= 2) begin: singleblock


memstream_singleblock
#(
    .CONFIG_EN(CONFIG_EN),
    .NSTREAMS(NSTREAMS),
    .MEM_DEPTH(MEM_DEPTH),
    .MEM_WIDTH(MEM_WIDTH),
    .MEM_INIT(MEM_INIT),
    .RAM_STYLE(RAM_STYLE),

    //widths per stream
    .STRM0_WIDTH(STRM0_WIDTH),
    .STRM1_WIDTH(STRM1_WIDTH),

    //depths per stream
    .STRM0_DEPTH(STRM0_DEPTH),
    .STRM1_DEPTH(STRM1_DEPTH),

    //offsets for each stream
    .STRM0_OFFSET(STRM0_OFFSET),
    .STRM1_OFFSET(STRM1_OFFSET)
)
mem
(
    .aclk(aclk),
    .aresetn(aresetn),

    .config_address(config_address),
    .config_ce(config_ce),
    .config_we(config_we),
    .config_d0(config_d0),
    .config_q0(config_q0),
    .config_rack(config_rack),

    .m_axis_0_tready(m_axis_0_tready),
    .m_axis_0_tvalid(m_axis_0_tvalid),
    .m_axis_0_tdata(m_axis_0_tdata),

    .m_axis_1_tready(m_axis_1_tready),
    .m_axis_1_tvalid(m_axis_1_tvalid),
    .m_axis_1_tdata(m_axis_1_tdata)
);

assign m_axis_2_tvalid = 0;
assign m_axis_2_tdata = 0;
assign m_axis_3_tvalid = 0;
assign m_axis_3_tdata = 0;
assign m_axis_4_tvalid = 0;
assign m_axis_4_tdata = 0;
assign m_axis_5_tvalid = 0;
assign m_axis_5_tdata = 0;

end else begin: multiblock


memstream_multiblock
#(
    .CONFIG_EN(CONFIG_EN),
    .NSTREAMS(NSTREAMS),
    .MEM_DEPTH(MEM_DEPTH),
    .MEM_WIDTH(MEM_WIDTH),
    .MEM_INIT(MEM_INIT),
    .RAM_STYLE(RAM_STYLE),

    //widths per stream
    .STRM0_WIDTH(STRM0_WIDTH),
    .STRM1_WIDTH(STRM1_WIDTH),
    .STRM2_WIDTH(STRM2_WIDTH),
    .STRM3_WIDTH(STRM3_WIDTH),
    .STRM4_WIDTH(STRM4_WIDTH),
    .STRM5_WIDTH(STRM5_WIDTH),

    //depths per stream
    .STRM0_DEPTH(STRM0_DEPTH),
    .STRM1_DEPTH(STRM1_DEPTH),
    .STRM2_DEPTH(STRM2_DEPTH),
    .STRM3_DEPTH(STRM3_DEPTH),
    .STRM4_DEPTH(STRM4_DEPTH),
    .STRM5_DEPTH(STRM5_DEPTH),

    //offsets for each stream
    .STRM0_OFFSET(STRM0_OFFSET),
    .STRM1_OFFSET(STRM1_OFFSET),
    .STRM2_OFFSET(STRM2_OFFSET),
    .STRM3_OFFSET(STRM3_OFFSET),
    .STRM4_OFFSET(STRM4_OFFSET),
    .STRM5_OFFSET(STRM5_OFFSET)
)
mem
(
    .aclk(aclk),
    .aresetn(aresetn),

    .config_address(config_address),
    .config_ce(config_ce),
    .config_we(config_we),
    .config_d0(config_d0),
    .config_q0(config_q0),

    .m_axis_0_afull(m_axis_0_afull),
    .m_axis_0_tready(m_axis_0_tready),
    .m_axis_0_tvalid(m_axis_0_tvalid),
    .m_axis_0_tdata(m_axis_0_tdata),

    .m_axis_1_afull(m_axis_1_afull),
    .m_axis_1_tready(m_axis_1_tready),
    .m_axis_1_tvalid(m_axis_1_tvalid),
    .m_axis_1_tdata(m_axis_1_tdata),

    .m_axis_2_afull(m_axis_2_afull),
    .m_axis_2_tready(m_axis_2_tready),
    .m_axis_2_tvalid(m_axis_2_tvalid),
    .m_axis_2_tdata(m_axis_2_tdata),

    .m_axis_3_afull(m_axis_3_afull),
    .m_axis_3_tready(m_axis_3_tready),
    .m_axis_3_tvalid(m_axis_3_tvalid),
    .m_axis_3_tdata(m_axis_3_tdata),

    .m_axis_4_afull(m_axis_4_afull),
    .m_axis_4_tready(m_axis_4_tready),
    .m_axis_4_tvalid(m_axis_4_tvalid),
    .m_axis_4_tdata(m_axis_4_tdata),

    .m_axis_5_afull(m_axis_5_afull),
    .m_axis_5_tready(m_axis_5_tready),
    .m_axis_5_tvalid(m_axis_5_tvalid),
    .m_axis_5_tdata(m_axis_5_tdata)

);


end
endgenerate

axi4lite_if
#(
    .ADDR_WIDTH(AXILITE_ADDR_WIDTH),
    .DATA_WIDTH(32),
    .IP_DATA_WIDTH(MEM_WIDTH)
)
config_if
(
    //system signals
    .aclk(aclk),
    .aresetn(aresetn),

    //Write channels
    //write address
    .awready(awready),
    .awvalid(awvalid),
    .awaddr(awaddr),
    .awprot(awprot),
    //write data
    .wready(wready),
    .wvalid(wvalid),
    .wdata(wdata),
    .wstrb(wstrb),
    //burst response
    .bready(bready),
    .bvalid(bvalid),
    .bresp(bresp),

    //Read channels
    //read address
    .arready(arready),
    .arvalid(arvalid),
    .araddr(araddr),
    .arprot(arprot),
    //read data
    .rready(rready),
    .rvalid(rvalid),
    .rresp(rresp),
    .rdata(rdata),

    //IP-side interface
    .ip_en(config_ce),
    .ip_wen(config_we),
    .ip_addr(config_address),
    .ip_wdata(config_d0),
    .ip_rack(config_rack),
    .ip_rdata(config_q0)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actcud.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actcud_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actcud_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actcud(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actcud_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actcud_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccud.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccud_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 2;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccud_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccud(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd2;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccud_rom Thresholding_Batch_0_Thresholding_Batccud_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActQgW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActQgW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActQgW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActQgW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActQgW_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActQgW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActMgi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActMgi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActMgi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActMgi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActMgi_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActMgi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActXh4.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActXh4_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActXh4_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActXh4(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActXh4_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActXh4_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/abe7/hdl/verilog/ConvolutionInputGenerator_0_ConvolutionInputGenerator_0.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="ConvolutionInputGenerator_0_ConvolutionInputGenerator_0,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=7.863750,HLS_SYN_LAT=59909,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=414,HLS_SYN_LUT=1768,HLS_VERSION=2020_1_1}" *)

module ConvolutionInputGenerator_0_ConvolutionInputGenerator_0 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [7:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_ConvolutionInputGene_1_fu_26_ap_start;
wire    grp_ConvolutionInputGene_1_fu_26_ap_done;
wire    grp_ConvolutionInputGene_1_fu_26_ap_idle;
wire    grp_ConvolutionInputGene_1_fu_26_ap_ready;
wire    grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY;
wire   [7:0] grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA;
wire    grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID;
wire    grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY;
reg    grp_ConvolutionInputGene_1_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [7:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_ConvolutionInputGene_1_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

ConvolutionInputGenerator_0_ConvolutionInputGene_1 grp_ConvolutionInputGene_1_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_ConvolutionInputGene_1_fu_26_ap_start),
    .ap_done(grp_ConvolutionInputGene_1_fu_26_ap_done),
    .ap_idle(grp_ConvolutionInputGene_1_fu_26_ap_idle),
    .ap_ready(grp_ConvolutionInputGene_1_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA),
    .vld_in(grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_ConvolutionInputGene_1_fu_26_ap_ready == 1'b1)) begin
            grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_ConvolutionInputGene_1_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_ConvolutionInputGene_1_fu_26_ap_start = grp_ConvolutionInputGene_1_fu_26_ap_start_reg;

assign grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //ConvolutionInputGenerator_0_ConvolutionInputGenerator_0
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc6D.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcc6D_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc6D_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcc6D(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcc6D_rom Thresholding_Batch_0_Thresholding_Batcc6D_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/b054/StreamingFIFO_14.v


module StreamingFIFO_14(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(16)
)
StreamingFIFO_14_StreamingFIFO_14
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/6c99/StreamingFIFO_8.v


module StreamingFIFO_8(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [31:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(32)
)
StreamingFIFO_8_StreamingFIFO_8
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccrw.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccrw_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccrw_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccrw(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccrw_rom Thresholding_Batch_0_Thresholding_Batccrw_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4c0f/hdl/verilog/StreamingDataWidthConverter_Batch_0_StreamingDataWidthConverter_Batch_0.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingDataWidthConverter_Batch_0_StreamingDataWidthConverter_Batch_0,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=5.025000,HLS_SYN_LAT=3077,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=95,HLS_SYN_LUT=213,HLS_VERSION=2020_1_1}" *)

module StreamingDataWidthConverter_Batch_0_StreamingDataWidthConverter_Batch_0 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [7:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [23:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_start;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_done;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_idle;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_ready;
wire    grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
wire   [23:0] grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY;
reg    grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [7:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_StreamingDataWidthCo_1_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingDataWidthConverter_Batch_0_StreamingDataWidthCo_1 grp_StreamingDataWidthCo_1_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_StreamingDataWidthCo_1_fu_26_ap_start),
    .ap_done(grp_StreamingDataWidthCo_1_fu_26_ap_done),
    .ap_idle(grp_StreamingDataWidthCo_1_fu_26_ap_idle),
    .ap_ready(grp_StreamingDataWidthCo_1_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 24 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .vld_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_StreamingDataWidthCo_1_fu_26_ap_ready == 1'b1)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_StreamingDataWidthCo_1_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_StreamingDataWidthCo_1_fu_26_ap_start = grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;

assign grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingDataWidthConverter_Batch_0_StreamingDataWidthConverter_Batch_0
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/2c22/hdl/verilog/ConvolutionInputGenerator_2_ConvolutionInputGene_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module ConvolutionInputGenerator_2_ConvolutionInputGene_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [23:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [23:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln197_fu_372_p2;
wire   [0:0] icmp_ln199_fu_394_p2;
wire   [0:0] and_ln245_fu_598_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln199_reg_885;
reg   [0:0] icmp_ln215_reg_889;
reg   [13:0] i_0_0_reg_275;
reg    ap_predicate_op117_read_state2;
reg    ap_predicate_op160_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_predicate_op203_write_state3;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [13:0] add_ln197_fu_378_p2;
wire   [0:0] icmp_ln215_fu_403_p2;
wire   [1:0] add_ln221_fu_461_p2;
reg   [1:0] add_ln221_reg_893;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
wire   [4:0] inputBuf_0_V_address0;
reg    inputBuf_0_V_ce0;
wire   [23:0] inputBuf_0_V_q0;
reg   [4:0] inputBuf_0_V_address1;
reg    inputBuf_0_V_ce1;
reg    inputBuf_0_V_we1;
wire   [4:0] inputBuf_1_V_address0;
reg    inputBuf_1_V_ce0;
wire   [23:0] inputBuf_1_V_q0;
reg   [4:0] inputBuf_1_V_address1;
reg    inputBuf_1_V_ce1;
reg    inputBuf_1_V_we1;
wire   [4:0] inputBuf_2_V_address0;
reg    inputBuf_2_V_ce0;
wire   [23:0] inputBuf_2_V_q0;
reg   [4:0] inputBuf_2_V_address1;
reg    inputBuf_2_V_ce1;
reg    inputBuf_2_V_we1;
wire   [4:0] inputBuf_3_V_address0;
reg    inputBuf_3_V_ce0;
wire   [23:0] inputBuf_3_V_q0;
reg   [4:0] inputBuf_3_V_address1;
reg    inputBuf_3_V_ce1;
reg    inputBuf_3_V_we1;
wire   [63:0] zext_ln221_fu_447_p1;
wire   [63:0] zext_ln248_fu_604_p1;
wire   [63:0] zext_ln202_fu_716_p1;
reg   [31:0] ofm_y_1_0_fu_82;
wire   [31:0] select_ln236_1_fu_555_p3;
wire   [0:0] icmp_ln224_fu_473_p2;
wire   [0:0] icmp_ln227_fu_490_p2;
wire   [0:0] icmp_ln230_fu_501_p2;
wire   [0:0] icmp_ln233_fu_521_p2;
reg   [31:0] ofm_x_1_0_fu_86;
wire   [31:0] add_ln232_fu_515_p2;
reg   [31:0] k_y_1_0_fu_90;
wire   [31:0] add_ln216_fu_425_p2;
reg   [31:0] inp_15_0_fu_94;
wire   [31:0] select_ln236_fu_547_p3;
wire   [31:0] add_ln204_fu_728_p2;
reg   [31:0] k_x_1_0_fu_98;
wire   [31:0] add_ln226_fu_484_p2;
reg   [31:0] count_simd_1_0_fu_102;
wire   [31:0] add_ln223_fu_467_p2;
reg   [31:0] read_block_1_0_fu_106;
wire   [31:0] zext_ln252_fu_669_p1;
wire   [31:0] add_ln211_fu_764_p2;
wire   [0:0] icmp_ln205_fu_346_p2;
reg   [31:0] current_block_write_s_fu_110;
wire   [31:0] select_ln252_fu_645_p3;
wire   [31:0] select_ln208_fu_756_p3;
reg   [31:0] current_line_1_0_fu_114;
wire   [31:0] select_ln252_1_fu_653_p3;
wire   [31:0] grp_fu_334_p2;
reg   [31:0] counter_internal_blo_fu_118;
wire   [31:0] select_ln264_fu_703_p3;
wire   [23:0] tmp_V_1_fu_780_p6;
reg    ap_block_pp0_stage0_01001;
wire   [1:0] trunc_ln321_1_fu_612_p1;
wire   [1:0] trunc_ln321_fu_724_p1;
wire   [31:0] add_ln220_fu_435_p2;
wire   [31:0] add_ln220_1_fu_441_p2;
wire   [1:0] trunc_ln216_1_fu_431_p1;
wire   [1:0] add_ln221_1_fu_455_p2;
wire   [1:0] trunc_ln216_fu_421_p1;
wire   [31:0] add_ln235_fu_535_p2;
wire   [0:0] icmp_ln236_fu_541_p2;
wire   [26:0] tmp_1_fu_582_p4;
wire   [0:0] icmp_ln245_fu_576_p2;
wire   [0:0] icmp_ln245_1_fu_592_p2;
wire   [5:0] trunc_ln197_fu_390_p1;
wire   [31:0] add_ln256_fu_625_p2;
wire   [0:0] icmp_ln257_fu_631_p2;
wire   [0:0] icmp_ln252_fu_340_p2;
wire   [31:0] select_ln257_fu_637_p3;
wire   [5:0] add_ln256_1_fu_619_p2;
wire   [5:0] select_ln252_2_fu_661_p3;
wire   [31:0] add_ln263_fu_691_p2;
wire   [0:0] icmp_ln264_fu_697_p2;
wire   [31:0] add_ln207_fu_744_p2;
wire   [0:0] icmp_ln208_fu_750_p2;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_block_pp0;
reg    ap_predicate_op125_store_state2;
reg    ap_enable_operation_125;
reg    ap_enable_state2_pp0_iter0_stage0;
reg    ap_predicate_op66_load_state2;
reg    ap_enable_operation_66;
reg    ap_predicate_op200_load_state3;
reg    ap_enable_operation_200;
reg    ap_enable_state3_pp0_iter1_stage0;
reg    ap_predicate_op168_store_state2;
reg    ap_enable_operation_168;
reg    ap_predicate_op127_store_state2;
reg    ap_enable_operation_127;
reg    ap_predicate_op64_load_state2;
reg    ap_enable_operation_64;
reg    ap_predicate_op199_load_state3;
reg    ap_enable_operation_199;
reg    ap_predicate_op170_store_state2;
reg    ap_enable_operation_170;
reg    ap_predicate_op129_store_state2;
reg    ap_enable_operation_129;
reg    ap_predicate_op62_load_state2;
reg    ap_enable_operation_62;
reg    ap_predicate_op198_load_state3;
reg    ap_enable_operation_198;
reg    ap_predicate_op172_store_state2;
reg    ap_enable_operation_172;
reg    ap_predicate_op131_store_state2;
reg    ap_enable_operation_131;
reg    ap_predicate_op68_load_state2;
reg    ap_enable_operation_68;
reg    ap_predicate_op201_load_state3;
reg    ap_enable_operation_201;
reg    ap_predicate_op174_store_state2;
reg    ap_enable_operation_174;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_654;
reg    ap_condition_230;
reg    ap_condition_660;
reg    ap_condition_664;
reg    ap_condition_668;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

ConvolutionInputGenerator_2_ConvolutionInputGbkb #(
    .DataWidth( 24 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
inputBuf_0_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_0_V_address0),
    .ce0(inputBuf_0_V_ce0),
    .q0(inputBuf_0_V_q0),
    .address1(inputBuf_0_V_address1),
    .ce1(inputBuf_0_V_ce1),
    .we1(inputBuf_0_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_2_ConvolutionInputGbkb #(
    .DataWidth( 24 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
inputBuf_1_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_1_V_address0),
    .ce0(inputBuf_1_V_ce0),
    .q0(inputBuf_1_V_q0),
    .address1(inputBuf_1_V_address1),
    .ce1(inputBuf_1_V_ce1),
    .we1(inputBuf_1_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_2_ConvolutionInputGbkb #(
    .DataWidth( 24 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
inputBuf_2_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_2_V_address0),
    .ce0(inputBuf_2_V_ce0),
    .q0(inputBuf_2_V_q0),
    .address1(inputBuf_2_V_address1),
    .ce1(inputBuf_2_V_ce1),
    .we1(inputBuf_2_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_2_ConvolutionInputGbkb #(
    .DataWidth( 24 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
inputBuf_3_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_3_V_address0),
    .ce0(inputBuf_3_V_ce0),
    .q0(inputBuf_3_V_q0),
    .address1(inputBuf_3_V_address1),
    .ce1(inputBuf_3_V_ce1),
    .we1(inputBuf_3_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_2_ConvolutionInputGfYi #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 24 ),
    .din1_WIDTH( 24 ),
    .din2_WIDTH( 24 ),
    .din3_WIDTH( 24 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 24 ))
ConvolutionInputGfYi_U1(
    .din0(inputBuf_0_V_q0),
    .din1(inputBuf_1_V_q0),
    .din2(inputBuf_2_V_q0),
    .din3(inputBuf_3_V_q0),
    .din4(add_ln221_reg_893),
    .dout(tmp_V_1_fu_780_p6)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln224_fu_473_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        count_simd_1_0_fu_102 <= add_ln223_fu_467_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln227_fu_490_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln230_fu_501_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln230_fu_501_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln233_fu_521_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln233_fu_521_p2 == 1'd1) & (icmp_ln230_fu_501_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        count_simd_1_0_fu_102 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        counter_internal_blo_fu_118 <= select_ln264_fu_703_p3;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_346_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        counter_internal_blo_fu_118 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_346_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_block_write_s_fu_110 <= select_ln208_fu_756_p3;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_block_write_s_fu_110 <= select_ln252_fu_645_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        current_block_write_s_fu_110 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln205_fu_346_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_line_1_0_fu_114 <= grp_fu_334_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_line_1_0_fu_114 <= select_ln252_1_fu_653_p3;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_346_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        current_line_1_0_fu_114 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_0_reg_275 <= 14'd0;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_0_reg_275 <= add_ln197_fu_378_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inp_15_0_fu_94 <= add_ln204_fu_728_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln233_fu_521_p2 == 1'd1) & (icmp_ln230_fu_501_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inp_15_0_fu_94 <= select_ln236_fu_547_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        inp_15_0_fu_94 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln227_fu_490_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        k_x_1_0_fu_98 <= add_ln226_fu_484_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln230_fu_501_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln230_fu_501_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln233_fu_521_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln233_fu_521_p2 == 1'd1) & (icmp_ln230_fu_501_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        k_x_1_0_fu_98 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln230_fu_501_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        k_y_1_0_fu_90 <= add_ln216_fu_425_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln230_fu_501_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        k_y_1_0_fu_90 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln230_fu_501_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln233_fu_521_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ofm_x_1_0_fu_86 <= add_ln232_fu_515_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln233_fu_521_p2 == 1'd1) & (icmp_ln230_fu_501_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ofm_x_1_0_fu_86 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln233_fu_521_p2 == 1'd1) & (icmp_ln230_fu_501_p2 == 1'd1) & (icmp_ln227_fu_490_p2 == 1'd1) & (icmp_ln224_fu_473_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ofm_y_1_0_fu_82 <= select_ln236_1_fu_555_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        ofm_y_1_0_fu_82 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_346_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        read_block_1_0_fu_106 <= add_ln211_fu_764_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        read_block_1_0_fu_106 <= zext_ln252_fu_669_p1;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        read_block_1_0_fu_106 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln221_reg_893 <= add_ln221_fu_461_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln197_fu_372_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln199_reg_885 <= icmp_ln199_fu_394_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln215_reg_889 <= icmp_ln215_fu_403_p2;
    end
end

always @ (*) begin
    if ((icmp_ln197_fu_372_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op160_read_state2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op117_read_state2 == 1'b1)))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_394_p2 == 1'd1) & (trunc_ln321_fu_724_p1 == 2'd0))) begin
            inputBuf_0_V_address1 = zext_ln202_fu_716_p1;
        end else if ((1'b1 == ap_condition_654)) begin
            inputBuf_0_V_address1 = zext_ln248_fu_604_p1;
        end else begin
            inputBuf_0_V_address1 = 'bx;
        end
    end else begin
        inputBuf_0_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_0_V_ce0 = 1'b1;
    end else begin
        inputBuf_0_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_0_V_ce1 = 1'b1;
    end else begin
        inputBuf_0_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_0_V_we1 = 1'b1;
    end else begin
        inputBuf_0_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_394_p2 == 1'd1) & (trunc_ln321_fu_724_p1 == 2'd1))) begin
            inputBuf_1_V_address1 = zext_ln202_fu_716_p1;
        end else if ((1'b1 == ap_condition_660)) begin
            inputBuf_1_V_address1 = zext_ln248_fu_604_p1;
        end else begin
            inputBuf_1_V_address1 = 'bx;
        end
    end else begin
        inputBuf_1_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_1_V_ce0 = 1'b1;
    end else begin
        inputBuf_1_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_1_V_ce1 = 1'b1;
    end else begin
        inputBuf_1_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_1_V_we1 = 1'b1;
    end else begin
        inputBuf_1_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_394_p2 == 1'd1) & (trunc_ln321_fu_724_p1 == 2'd2))) begin
            inputBuf_2_V_address1 = zext_ln202_fu_716_p1;
        end else if ((1'b1 == ap_condition_664)) begin
            inputBuf_2_V_address1 = zext_ln248_fu_604_p1;
        end else begin
            inputBuf_2_V_address1 = 'bx;
        end
    end else begin
        inputBuf_2_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_2_V_ce0 = 1'b1;
    end else begin
        inputBuf_2_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_2_V_ce1 = 1'b1;
    end else begin
        inputBuf_2_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_2_V_we1 = 1'b1;
    end else begin
        inputBuf_2_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_394_p2 == 1'd1) & (trunc_ln321_fu_724_p1 == 2'd3))) begin
            inputBuf_3_V_address1 = zext_ln202_fu_716_p1;
        end else if ((1'b1 == ap_condition_668)) begin
            inputBuf_3_V_address1 = zext_ln248_fu_604_p1;
        end else begin
            inputBuf_3_V_address1 = 'bx;
        end
    end else begin
        inputBuf_3_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_3_V_ce0 = 1'b1;
    end else begin
        inputBuf_3_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_3_V_ce1 = 1'b1;
    end else begin
        inputBuf_3_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_3_V_we1 = 1'b1;
    end else begin
        inputBuf_3_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln215_reg_889 == 1'd1) & (icmp_ln199_reg_885 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op203_write_state3 == 1'b1))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((icmp_ln197_fu_372_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((icmp_ln197_fu_372_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln197_fu_378_p2 = (i_0_0_reg_275 + 14'd1);

assign add_ln204_fu_728_p2 = (inp_15_0_fu_94 + 32'd1);

assign add_ln207_fu_744_p2 = (current_block_write_s_fu_110 + 32'd1);

assign add_ln211_fu_764_p2 = (read_block_1_0_fu_106 + 32'd1);

assign add_ln216_fu_425_p2 = (32'd1 + k_y_1_0_fu_90);

assign add_ln220_1_fu_441_p2 = (add_ln220_fu_435_p2 + k_x_1_0_fu_98);

assign add_ln220_fu_435_p2 = (ofm_x_1_0_fu_86 + count_simd_1_0_fu_102);

assign add_ln221_1_fu_455_p2 = (2'd1 + trunc_ln216_1_fu_431_p1);

assign add_ln221_fu_461_p2 = (add_ln221_1_fu_455_p2 + trunc_ln216_fu_421_p1);

assign add_ln223_fu_467_p2 = (32'd1 + count_simd_1_0_fu_102);

assign add_ln226_fu_484_p2 = (k_x_1_0_fu_98 + 32'd1);

assign add_ln232_fu_515_p2 = (ofm_x_1_0_fu_86 + 32'd1);

assign add_ln235_fu_535_p2 = (ofm_y_1_0_fu_82 + 32'd1);

assign add_ln256_1_fu_619_p2 = (trunc_ln197_fu_390_p1 + 6'd1);

assign add_ln256_fu_625_p2 = (current_block_write_s_fu_110 + 32'd1);

assign add_ln263_fu_691_p2 = (counter_internal_blo_fu_118 + 32'd1);

assign and_ln245_fu_598_p2 = (icmp_ln245_fu_576_p2 & icmp_ln245_1_fu_592_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

always @ (*) begin
    ap_block_pp0 = ((ap_ST_fsm_pp0_stage0 == ap_CS_fsm) & (1'b1 == ap_block_pp0_stage0_subdone));
end

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op160_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op117_read_state2 == 1'b1))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op160_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op117_read_state2 == 1'b1)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op160_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op117_read_state2 == 1'b1)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op160_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op117_read_state2 == 1'b1)));
end

always @ (*) begin
    ap_block_state3_io = ((out_V_V_TREADY == 1'b0) & (ap_predicate_op203_write_state3 == 1'b1));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_230 = ((icmp_ln197_fu_372_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_condition_654 = ((1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd0));
end

always @ (*) begin
    ap_condition_660 = ((1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd1));
end

always @ (*) begin
    ap_condition_664 = ((1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd2));
end

always @ (*) begin
    ap_condition_668 = ((1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd3));
end

always @ (*) begin
    ap_enable_operation_125 = (ap_predicate_op125_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_127 = (ap_predicate_op127_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_129 = (ap_predicate_op129_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_131 = (ap_predicate_op131_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_168 = (ap_predicate_op168_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_170 = (ap_predicate_op170_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_172 = (ap_predicate_op172_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_174 = (ap_predicate_op174_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_198 = (ap_predicate_op198_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_199 = (ap_predicate_op199_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_200 = (ap_predicate_op200_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_201 = (ap_predicate_op201_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_62 = (ap_predicate_op62_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_64 = (ap_predicate_op64_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_66 = (ap_predicate_op66_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_68 = (ap_predicate_op68_load_state2 == 1'b1);
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

always @ (*) begin
    ap_enable_state2_pp0_iter0_stage0 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_enable_state3_pp0_iter1_stage0 = ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_predicate_op117_read_state2 = ((1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op125_store_state2 = ((1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd2));
end

always @ (*) begin
    ap_predicate_op127_store_state2 = ((1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd1));
end

always @ (*) begin
    ap_predicate_op129_store_state2 = ((1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd0));
end

always @ (*) begin
    ap_predicate_op131_store_state2 = ((1'd1 == and_ln245_fu_598_p2) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_1_fu_612_p1 == 2'd3));
end

always @ (*) begin
    ap_predicate_op160_read_state2 = ((icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op168_store_state2 = ((icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd2));
end

always @ (*) begin
    ap_predicate_op170_store_state2 = ((icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd1));
end

always @ (*) begin
    ap_predicate_op172_store_state2 = ((icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd0));
end

always @ (*) begin
    ap_predicate_op174_store_state2 = ((icmp_ln199_fu_394_p2 == 1'd1) & (icmp_ln197_fu_372_p2 == 1'd0) & (trunc_ln321_fu_724_p1 == 2'd3));
end

always @ (*) begin
    ap_predicate_op198_load_state3 = ((icmp_ln215_reg_889 == 1'd1) & (icmp_ln199_reg_885 == 1'd0));
end

always @ (*) begin
    ap_predicate_op199_load_state3 = ((icmp_ln215_reg_889 == 1'd1) & (icmp_ln199_reg_885 == 1'd0));
end

always @ (*) begin
    ap_predicate_op200_load_state3 = ((icmp_ln215_reg_889 == 1'd1) & (icmp_ln199_reg_885 == 1'd0));
end

always @ (*) begin
    ap_predicate_op201_load_state3 = ((icmp_ln215_reg_889 == 1'd1) & (icmp_ln199_reg_885 == 1'd0));
end

always @ (*) begin
    ap_predicate_op203_write_state3 = ((icmp_ln215_reg_889 == 1'd1) & (icmp_ln199_reg_885 == 1'd0));
end

always @ (*) begin
    ap_predicate_op62_load_state2 = ((icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op64_load_state2 = ((icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op66_load_state2 = ((icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op68_load_state2 = ((icmp_ln215_fu_403_p2 == 1'd1) & (icmp_ln199_fu_394_p2 == 1'd0) & (icmp_ln197_fu_372_p2 == 1'd0));
end

assign grp_fu_334_p2 = (current_line_1_0_fu_114 + 32'd1);

assign icmp_ln197_fu_372_p2 = ((i_0_0_reg_275 == 14'd8196) ? 1'b1 : 1'b0);

assign icmp_ln199_fu_394_p2 = ((inp_15_0_fu_94 < 32'd96) ? 1'b1 : 1'b0);

assign icmp_ln205_fu_346_p2 = ((grp_fu_334_p2 == 32'd32) ? 1'b1 : 1'b0);

assign icmp_ln208_fu_750_p2 = ((add_ln207_fu_744_p2 == 32'd4) ? 1'b1 : 1'b0);

assign icmp_ln215_fu_403_p2 = ((counter_internal_blo_fu_118 < 32'd269) ? 1'b1 : 1'b0);

assign icmp_ln224_fu_473_p2 = ((count_simd_1_0_fu_102 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln227_fu_490_p2 = ((add_ln226_fu_484_p2 == 32'd3) ? 1'b1 : 1'b0);

assign icmp_ln230_fu_501_p2 = ((add_ln216_fu_425_p2 == 32'd3) ? 1'b1 : 1'b0);

assign icmp_ln233_fu_521_p2 = ((add_ln232_fu_515_p2 == 32'd30) ? 1'b1 : 1'b0);

assign icmp_ln236_fu_541_p2 = ((add_ln235_fu_535_p2 == 32'd30) ? 1'b1 : 1'b0);

assign icmp_ln245_1_fu_592_p2 = ((tmp_1_fu_582_p4 == 27'd0) ? 1'b1 : 1'b0);

assign icmp_ln245_fu_576_p2 = ((counter_internal_blo_fu_118 < 32'd31) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_340_p2 = ((grp_fu_334_p2 == 32'd32) ? 1'b1 : 1'b0);

assign icmp_ln257_fu_631_p2 = ((add_ln256_fu_625_p2 == 32'd4) ? 1'b1 : 1'b0);

assign icmp_ln264_fu_697_p2 = ((add_ln263_fu_691_p2 == 32'd269) ? 1'b1 : 1'b0);

assign inputBuf_0_V_address0 = zext_ln221_fu_447_p1;

assign inputBuf_1_V_address0 = zext_ln221_fu_447_p1;

assign inputBuf_2_V_address0 = zext_ln221_fu_447_p1;

assign inputBuf_3_V_address0 = zext_ln221_fu_447_p1;

assign out_V_V_TDATA = tmp_V_1_fu_780_p6;

assign select_ln208_fu_756_p3 = ((icmp_ln208_fu_750_p2[0:0] === 1'b1) ? 32'd0 : add_ln207_fu_744_p2);

assign select_ln236_1_fu_555_p3 = ((icmp_ln236_fu_541_p2[0:0] === 1'b1) ? 32'd0 : add_ln235_fu_535_p2);

assign select_ln236_fu_547_p3 = ((icmp_ln236_fu_541_p2[0:0] === 1'b1) ? 32'd0 : inp_15_0_fu_94);

assign select_ln252_1_fu_653_p3 = ((icmp_ln252_fu_340_p2[0:0] === 1'b1) ? 32'd0 : grp_fu_334_p2);

assign select_ln252_2_fu_661_p3 = ((icmp_ln252_fu_340_p2[0:0] === 1'b1) ? add_ln256_1_fu_619_p2 : trunc_ln197_fu_390_p1);

assign select_ln252_fu_645_p3 = ((icmp_ln252_fu_340_p2[0:0] === 1'b1) ? select_ln257_fu_637_p3 : current_block_write_s_fu_110);

assign select_ln257_fu_637_p3 = ((icmp_ln257_fu_631_p2[0:0] === 1'b1) ? 32'd0 : add_ln256_fu_625_p2);

assign select_ln264_fu_703_p3 = ((icmp_ln264_fu_697_p2[0:0] === 1'b1) ? 32'd0 : add_ln263_fu_691_p2);

assign tmp_1_fu_582_p4 = {{read_block_1_0_fu_106[31:5]}};

assign trunc_ln197_fu_390_p1 = read_block_1_0_fu_106[5:0];

assign trunc_ln216_1_fu_431_p1 = current_block_write_s_fu_110[1:0];

assign trunc_ln216_fu_421_p1 = k_y_1_0_fu_90[1:0];

assign trunc_ln321_1_fu_612_p1 = current_block_write_s_fu_110[1:0];

assign trunc_ln321_fu_724_p1 = current_block_write_s_fu_110[1:0];

assign zext_ln202_fu_716_p1 = current_line_1_0_fu_114;

assign zext_ln221_fu_447_p1 = add_ln220_1_fu_441_p2;

assign zext_ln248_fu_604_p1 = current_line_1_0_fu_114;

assign zext_ln252_fu_669_p1 = select_ln252_2_fu_661_p3;

endmodule //ConvolutionInputGenerator_2_ConvolutionInputGene_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccEy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccEy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccEy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccEy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccEy_rom Thresholding_Batch_0_Thresholding_BatccEy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_StreamingFCLayer_5jm.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module StreamingFCLayer_Batch_1_StreamingFCLayer_5jm #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH       = 32,
    din5_WIDTH       = 32,
    din6_WIDTH       = 32,
    din7_WIDTH       = 32,
    din8_WIDTH       = 32,
    din9_WIDTH       = 32,
    din10_WIDTH       = 32,
    din11_WIDTH       = 32,
    din12_WIDTH       = 32,
    din13_WIDTH       = 32,
    din14_WIDTH       = 32,
    din15_WIDTH       = 32,
    din16_WIDTH       = 32,
    din17_WIDTH       = 32,
    din18_WIDTH       = 32,
    din19_WIDTH       = 32,
    din20_WIDTH       = 32,
    din21_WIDTH       = 32,
    din22_WIDTH       = 32,
    din23_WIDTH       = 32,
    din24_WIDTH       = 32,
    din25_WIDTH       = 32,
    din26_WIDTH       = 32,
    din27_WIDTH       = 32,
    din28_WIDTH       = 32,
    din29_WIDTH       = 32,
    din30_WIDTH       = 32,
    din31_WIDTH       = 32,
    din32_WIDTH       = 32,
    din33_WIDTH       = 32,
    din34_WIDTH       = 32,
    din35_WIDTH       = 32,
    din36_WIDTH       = 32,
    din37_WIDTH       = 32,
    din38_WIDTH       = 32,
    din39_WIDTH       = 32,
    din40_WIDTH       = 32,
    din41_WIDTH       = 32,
    din42_WIDTH       = 32,
    din43_WIDTH       = 32,
    din44_WIDTH       = 32,
    din45_WIDTH       = 32,
    din46_WIDTH       = 32,
    din47_WIDTH       = 32,
    din48_WIDTH       = 32,
    din49_WIDTH       = 32,
    din50_WIDTH       = 32,
    din51_WIDTH       = 32,
    din52_WIDTH       = 32,
    din53_WIDTH       = 32,
    din54_WIDTH       = 32,
    din55_WIDTH       = 32,
    din56_WIDTH       = 32,
    din57_WIDTH       = 32,
    din58_WIDTH       = 32,
    din59_WIDTH       = 32,
    din60_WIDTH       = 32,
    din61_WIDTH       = 32,
    din62_WIDTH       = 32,
    din63_WIDTH       = 32,
    din64_WIDTH       = 32,
    din65_WIDTH       = 32,
    din66_WIDTH       = 32,
    din67_WIDTH       = 32,
    din68_WIDTH       = 32,
    din69_WIDTH       = 32,
    din70_WIDTH       = 32,
    din71_WIDTH       = 32,
    din72_WIDTH       = 32,
    din73_WIDTH       = 32,
    din74_WIDTH       = 32,
    din75_WIDTH       = 32,
    din76_WIDTH       = 32,
    din77_WIDTH       = 32,
    din78_WIDTH       = 32,
    din79_WIDTH       = 32,
    din80_WIDTH       = 32,
    din81_WIDTH       = 32,
    din82_WIDTH       = 32,
    din83_WIDTH       = 32,
    din84_WIDTH       = 32,
    din85_WIDTH       = 32,
    din86_WIDTH       = 32,
    din87_WIDTH       = 32,
    din88_WIDTH       = 32,
    din89_WIDTH       = 32,
    din90_WIDTH       = 32,
    din91_WIDTH       = 32,
    din92_WIDTH       = 32,
    din93_WIDTH       = 32,
    din94_WIDTH       = 32,
    din95_WIDTH       = 32,
    din96_WIDTH       = 32,
    din97_WIDTH       = 32,
    din98_WIDTH       = 32,
    din99_WIDTH       = 32,
    din100_WIDTH       = 32,
    din101_WIDTH       = 32,
    din102_WIDTH       = 32,
    din103_WIDTH       = 32,
    din104_WIDTH       = 32,
    din105_WIDTH       = 32,
    din106_WIDTH       = 32,
    din107_WIDTH       = 32,
    din108_WIDTH       = 32,
    din109_WIDTH       = 32,
    din110_WIDTH       = 32,
    din111_WIDTH       = 32,
    din112_WIDTH       = 32,
    din113_WIDTH       = 32,
    din114_WIDTH       = 32,
    din115_WIDTH       = 32,
    din116_WIDTH       = 32,
    din117_WIDTH       = 32,
    din118_WIDTH       = 32,
    din119_WIDTH       = 32,
    din120_WIDTH       = 32,
    din121_WIDTH       = 32,
    din122_WIDTH       = 32,
    din123_WIDTH       = 32,
    din124_WIDTH       = 32,
    din125_WIDTH       = 32,
    din126_WIDTH       = 32,
    din127_WIDTH       = 32,
    din128_WIDTH       = 32,
    din129_WIDTH       = 32,
    din130_WIDTH       = 32,
    din131_WIDTH       = 32,
    din132_WIDTH       = 32,
    din133_WIDTH       = 32,
    din134_WIDTH       = 32,
    din135_WIDTH       = 32,
    din136_WIDTH       = 32,
    din137_WIDTH       = 32,
    din138_WIDTH       = 32,
    din139_WIDTH       = 32,
    din140_WIDTH       = 32,
    din141_WIDTH       = 32,
    din142_WIDTH       = 32,
    din143_WIDTH       = 32,
    din144_WIDTH       = 32,
    din145_WIDTH       = 32,
    din146_WIDTH       = 32,
    din147_WIDTH       = 32,
    din148_WIDTH       = 32,
    din149_WIDTH       = 32,
    din150_WIDTH       = 32,
    din151_WIDTH       = 32,
    din152_WIDTH       = 32,
    din153_WIDTH       = 32,
    din154_WIDTH       = 32,
    din155_WIDTH       = 32,
    din156_WIDTH       = 32,
    din157_WIDTH       = 32,
    din158_WIDTH       = 32,
    din159_WIDTH       = 32,
    din160_WIDTH       = 32,
    din161_WIDTH       = 32,
    din162_WIDTH       = 32,
    din163_WIDTH       = 32,
    din164_WIDTH       = 32,
    din165_WIDTH       = 32,
    din166_WIDTH       = 32,
    din167_WIDTH       = 32,
    din168_WIDTH       = 32,
    din169_WIDTH       = 32,
    din170_WIDTH       = 32,
    din171_WIDTH       = 32,
    din172_WIDTH       = 32,
    din173_WIDTH       = 32,
    din174_WIDTH       = 32,
    din175_WIDTH       = 32,
    din176_WIDTH       = 32,
    din177_WIDTH       = 32,
    din178_WIDTH       = 32,
    din179_WIDTH       = 32,
    din180_WIDTH       = 32,
    din181_WIDTH       = 32,
    din182_WIDTH       = 32,
    din183_WIDTH       = 32,
    din184_WIDTH       = 32,
    din185_WIDTH       = 32,
    din186_WIDTH       = 32,
    din187_WIDTH       = 32,
    din188_WIDTH       = 32,
    din189_WIDTH       = 32,
    din190_WIDTH       = 32,
    din191_WIDTH       = 32,
    din192_WIDTH       = 32,
    din193_WIDTH       = 32,
    din194_WIDTH       = 32,
    din195_WIDTH       = 32,
    din196_WIDTH       = 32,
    din197_WIDTH       = 32,
    din198_WIDTH       = 32,
    din199_WIDTH       = 32,
    din200_WIDTH       = 32,
    din201_WIDTH       = 32,
    din202_WIDTH       = 32,
    din203_WIDTH       = 32,
    din204_WIDTH       = 32,
    din205_WIDTH       = 32,
    din206_WIDTH       = 32,
    din207_WIDTH       = 32,
    din208_WIDTH       = 32,
    din209_WIDTH       = 32,
    din210_WIDTH       = 32,
    din211_WIDTH       = 32,
    din212_WIDTH       = 32,
    din213_WIDTH       = 32,
    din214_WIDTH       = 32,
    din215_WIDTH       = 32,
    din216_WIDTH       = 32,
    din217_WIDTH       = 32,
    din218_WIDTH       = 32,
    din219_WIDTH       = 32,
    din220_WIDTH       = 32,
    din221_WIDTH       = 32,
    din222_WIDTH       = 32,
    din223_WIDTH       = 32,
    din224_WIDTH       = 32,
    din225_WIDTH       = 32,
    din226_WIDTH       = 32,
    din227_WIDTH       = 32,
    din228_WIDTH       = 32,
    din229_WIDTH       = 32,
    din230_WIDTH       = 32,
    din231_WIDTH       = 32,
    din232_WIDTH       = 32,
    din233_WIDTH       = 32,
    din234_WIDTH       = 32,
    din235_WIDTH       = 32,
    din236_WIDTH       = 32,
    din237_WIDTH       = 32,
    din238_WIDTH       = 32,
    din239_WIDTH       = 32,
    din240_WIDTH       = 32,
    din241_WIDTH       = 32,
    din242_WIDTH       = 32,
    din243_WIDTH       = 32,
    din244_WIDTH       = 32,
    din245_WIDTH       = 32,
    din246_WIDTH       = 32,
    din247_WIDTH       = 32,
    din248_WIDTH       = 32,
    din249_WIDTH       = 32,
    din250_WIDTH       = 32,
    din251_WIDTH       = 32,
    din252_WIDTH       = 32,
    din253_WIDTH       = 32,
    din254_WIDTH       = 32,
    din255_WIDTH       = 32,
    din256_WIDTH       = 32,
    din257_WIDTH       = 32,
    din258_WIDTH       = 32,
    din259_WIDTH       = 32,
    din260_WIDTH       = 32,
    din261_WIDTH       = 32,
    din262_WIDTH       = 32,
    din263_WIDTH       = 32,
    din264_WIDTH       = 32,
    din265_WIDTH       = 32,
    din266_WIDTH       = 32,
    din267_WIDTH       = 32,
    din268_WIDTH       = 32,
    din269_WIDTH       = 32,
    din270_WIDTH       = 32,
    din271_WIDTH       = 32,
    din272_WIDTH       = 32,
    din273_WIDTH       = 32,
    din274_WIDTH       = 32,
    din275_WIDTH       = 32,
    din276_WIDTH       = 32,
    din277_WIDTH       = 32,
    din278_WIDTH       = 32,
    din279_WIDTH       = 32,
    din280_WIDTH       = 32,
    din281_WIDTH       = 32,
    din282_WIDTH       = 32,
    din283_WIDTH       = 32,
    din284_WIDTH       = 32,
    din285_WIDTH       = 32,
    din286_WIDTH       = 32,
    din287_WIDTH       = 32,
    din288_WIDTH       = 32,
    din289_WIDTH       = 32,
    din290_WIDTH       = 32,
    din291_WIDTH       = 32,
    din292_WIDTH       = 32,
    din293_WIDTH       = 32,
    din294_WIDTH       = 32,
    din295_WIDTH       = 32,
    din296_WIDTH       = 32,
    din297_WIDTH       = 32,
    din298_WIDTH       = 32,
    din299_WIDTH       = 32,
    din300_WIDTH       = 32,
    din301_WIDTH       = 32,
    din302_WIDTH       = 32,
    din303_WIDTH       = 32,
    din304_WIDTH       = 32,
    din305_WIDTH       = 32,
    din306_WIDTH       = 32,
    din307_WIDTH       = 32,
    din308_WIDTH       = 32,
    din309_WIDTH       = 32,
    din310_WIDTH       = 32,
    din311_WIDTH       = 32,
    din312_WIDTH       = 32,
    din313_WIDTH       = 32,
    din314_WIDTH       = 32,
    din315_WIDTH       = 32,
    din316_WIDTH       = 32,
    din317_WIDTH       = 32,
    din318_WIDTH       = 32,
    din319_WIDTH       = 32,
    din320_WIDTH       = 32,
    din321_WIDTH       = 32,
    din322_WIDTH       = 32,
    din323_WIDTH       = 32,
    din324_WIDTH       = 32,
    din325_WIDTH       = 32,
    din326_WIDTH       = 32,
    din327_WIDTH       = 32,
    din328_WIDTH       = 32,
    din329_WIDTH       = 32,
    din330_WIDTH       = 32,
    din331_WIDTH       = 32,
    din332_WIDTH       = 32,
    din333_WIDTH       = 32,
    din334_WIDTH       = 32,
    din335_WIDTH       = 32,
    din336_WIDTH       = 32,
    din337_WIDTH       = 32,
    din338_WIDTH       = 32,
    din339_WIDTH       = 32,
    din340_WIDTH       = 32,
    din341_WIDTH       = 32,
    din342_WIDTH       = 32,
    din343_WIDTH       = 32,
    din344_WIDTH       = 32,
    din345_WIDTH       = 32,
    din346_WIDTH       = 32,
    din347_WIDTH       = 32,
    din348_WIDTH       = 32,
    din349_WIDTH       = 32,
    din350_WIDTH       = 32,
    din351_WIDTH       = 32,
    din352_WIDTH       = 32,
    din353_WIDTH       = 32,
    din354_WIDTH       = 32,
    din355_WIDTH       = 32,
    din356_WIDTH       = 32,
    din357_WIDTH       = 32,
    din358_WIDTH       = 32,
    din359_WIDTH       = 32,
    din360_WIDTH       = 32,
    din361_WIDTH       = 32,
    din362_WIDTH       = 32,
    din363_WIDTH       = 32,
    din364_WIDTH       = 32,
    din365_WIDTH       = 32,
    din366_WIDTH       = 32,
    din367_WIDTH       = 32,
    din368_WIDTH       = 32,
    din369_WIDTH       = 32,
    din370_WIDTH       = 32,
    din371_WIDTH       = 32,
    din372_WIDTH       = 32,
    din373_WIDTH       = 32,
    din374_WIDTH       = 32,
    din375_WIDTH       = 32,
    din376_WIDTH       = 32,
    din377_WIDTH       = 32,
    din378_WIDTH       = 32,
    din379_WIDTH       = 32,
    din380_WIDTH       = 32,
    din381_WIDTH       = 32,
    din382_WIDTH       = 32,
    din383_WIDTH       = 32,
    din384_WIDTH       = 32,
    din385_WIDTH       = 32,
    din386_WIDTH       = 32,
    din387_WIDTH       = 32,
    din388_WIDTH       = 32,
    din389_WIDTH       = 32,
    din390_WIDTH       = 32,
    din391_WIDTH       = 32,
    din392_WIDTH       = 32,
    din393_WIDTH       = 32,
    din394_WIDTH       = 32,
    din395_WIDTH       = 32,
    din396_WIDTH       = 32,
    din397_WIDTH       = 32,
    din398_WIDTH       = 32,
    din399_WIDTH       = 32,
    din400_WIDTH       = 32,
    din401_WIDTH       = 32,
    din402_WIDTH       = 32,
    din403_WIDTH       = 32,
    din404_WIDTH       = 32,
    din405_WIDTH       = 32,
    din406_WIDTH       = 32,
    din407_WIDTH       = 32,
    din408_WIDTH       = 32,
    din409_WIDTH       = 32,
    din410_WIDTH       = 32,
    din411_WIDTH       = 32,
    din412_WIDTH       = 32,
    din413_WIDTH       = 32,
    din414_WIDTH       = 32,
    din415_WIDTH       = 32,
    din416_WIDTH       = 32,
    din417_WIDTH       = 32,
    din418_WIDTH       = 32,
    din419_WIDTH       = 32,
    din420_WIDTH       = 32,
    din421_WIDTH       = 32,
    din422_WIDTH       = 32,
    din423_WIDTH       = 32,
    din424_WIDTH       = 32,
    din425_WIDTH       = 32,
    din426_WIDTH       = 32,
    din427_WIDTH       = 32,
    din428_WIDTH       = 32,
    din429_WIDTH       = 32,
    din430_WIDTH       = 32,
    din431_WIDTH       = 32,
    din432_WIDTH       = 32,
    din433_WIDTH       = 32,
    din434_WIDTH       = 32,
    din435_WIDTH       = 32,
    din436_WIDTH       = 32,
    din437_WIDTH       = 32,
    din438_WIDTH       = 32,
    din439_WIDTH       = 32,
    din440_WIDTH       = 32,
    din441_WIDTH       = 32,
    din442_WIDTH       = 32,
    din443_WIDTH       = 32,
    din444_WIDTH       = 32,
    din445_WIDTH       = 32,
    din446_WIDTH       = 32,
    din447_WIDTH       = 32,
    din448_WIDTH       = 32,
    din449_WIDTH       = 32,
    din450_WIDTH       = 32,
    din451_WIDTH       = 32,
    din452_WIDTH       = 32,
    din453_WIDTH       = 32,
    din454_WIDTH       = 32,
    din455_WIDTH       = 32,
    din456_WIDTH       = 32,
    din457_WIDTH       = 32,
    din458_WIDTH       = 32,
    din459_WIDTH       = 32,
    din460_WIDTH       = 32,
    din461_WIDTH       = 32,
    din462_WIDTH       = 32,
    din463_WIDTH       = 32,
    din464_WIDTH       = 32,
    din465_WIDTH       = 32,
    din466_WIDTH       = 32,
    din467_WIDTH       = 32,
    din468_WIDTH       = 32,
    din469_WIDTH       = 32,
    din470_WIDTH       = 32,
    din471_WIDTH       = 32,
    din472_WIDTH       = 32,
    din473_WIDTH       = 32,
    din474_WIDTH       = 32,
    din475_WIDTH       = 32,
    din476_WIDTH       = 32,
    din477_WIDTH       = 32,
    din478_WIDTH       = 32,
    din479_WIDTH       = 32,
    din480_WIDTH       = 32,
    din481_WIDTH       = 32,
    din482_WIDTH       = 32,
    din483_WIDTH       = 32,
    din484_WIDTH       = 32,
    din485_WIDTH       = 32,
    din486_WIDTH       = 32,
    din487_WIDTH       = 32,
    din488_WIDTH       = 32,
    din489_WIDTH       = 32,
    din490_WIDTH       = 32,
    din491_WIDTH       = 32,
    din492_WIDTH       = 32,
    din493_WIDTH       = 32,
    din494_WIDTH       = 32,
    din495_WIDTH       = 32,
    din496_WIDTH       = 32,
    din497_WIDTH       = 32,
    din498_WIDTH       = 32,
    din499_WIDTH       = 32,
    din500_WIDTH       = 32,
    din501_WIDTH       = 32,
    din502_WIDTH       = 32,
    din503_WIDTH       = 32,
    din504_WIDTH       = 32,
    din505_WIDTH       = 32,
    din506_WIDTH       = 32,
    din507_WIDTH       = 32,
    din508_WIDTH       = 32,
    din509_WIDTH       = 32,
    din510_WIDTH       = 32,
    din511_WIDTH       = 32,
    din512_WIDTH       = 32,
    din513_WIDTH       = 32,
    din514_WIDTH       = 32,
    din515_WIDTH       = 32,
    din516_WIDTH       = 32,
    din517_WIDTH       = 32,
    din518_WIDTH       = 32,
    din519_WIDTH       = 32,
    din520_WIDTH       = 32,
    din521_WIDTH       = 32,
    din522_WIDTH       = 32,
    din523_WIDTH       = 32,
    din524_WIDTH       = 32,
    din525_WIDTH       = 32,
    din526_WIDTH       = 32,
    din527_WIDTH       = 32,
    din528_WIDTH       = 32,
    din529_WIDTH       = 32,
    din530_WIDTH       = 32,
    din531_WIDTH       = 32,
    din532_WIDTH       = 32,
    din533_WIDTH       = 32,
    din534_WIDTH       = 32,
    din535_WIDTH       = 32,
    din536_WIDTH       = 32,
    din537_WIDTH       = 32,
    din538_WIDTH       = 32,
    din539_WIDTH       = 32,
    din540_WIDTH       = 32,
    din541_WIDTH       = 32,
    din542_WIDTH       = 32,
    din543_WIDTH       = 32,
    din544_WIDTH       = 32,
    din545_WIDTH       = 32,
    din546_WIDTH       = 32,
    din547_WIDTH       = 32,
    din548_WIDTH       = 32,
    din549_WIDTH       = 32,
    din550_WIDTH       = 32,
    din551_WIDTH       = 32,
    din552_WIDTH       = 32,
    din553_WIDTH       = 32,
    din554_WIDTH       = 32,
    din555_WIDTH       = 32,
    din556_WIDTH       = 32,
    din557_WIDTH       = 32,
    din558_WIDTH       = 32,
    din559_WIDTH       = 32,
    din560_WIDTH       = 32,
    din561_WIDTH       = 32,
    din562_WIDTH       = 32,
    din563_WIDTH       = 32,
    din564_WIDTH       = 32,
    din565_WIDTH       = 32,
    din566_WIDTH       = 32,
    din567_WIDTH       = 32,
    din568_WIDTH       = 32,
    din569_WIDTH       = 32,
    din570_WIDTH       = 32,
    din571_WIDTH       = 32,
    din572_WIDTH       = 32,
    din573_WIDTH       = 32,
    din574_WIDTH       = 32,
    din575_WIDTH       = 32,
    din576_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [15 : 0]     din0,
    input  [15 : 0]     din1,
    input  [15 : 0]     din2,
    input  [15 : 0]     din3,
    input  [15 : 0]     din4,
    input  [15 : 0]     din5,
    input  [15 : 0]     din6,
    input  [15 : 0]     din7,
    input  [15 : 0]     din8,
    input  [15 : 0]     din9,
    input  [15 : 0]     din10,
    input  [15 : 0]     din11,
    input  [15 : 0]     din12,
    input  [15 : 0]     din13,
    input  [15 : 0]     din14,
    input  [15 : 0]     din15,
    input  [15 : 0]     din16,
    input  [15 : 0]     din17,
    input  [15 : 0]     din18,
    input  [15 : 0]     din19,
    input  [15 : 0]     din20,
    input  [15 : 0]     din21,
    input  [15 : 0]     din22,
    input  [15 : 0]     din23,
    input  [15 : 0]     din24,
    input  [15 : 0]     din25,
    input  [15 : 0]     din26,
    input  [15 : 0]     din27,
    input  [15 : 0]     din28,
    input  [15 : 0]     din29,
    input  [15 : 0]     din30,
    input  [15 : 0]     din31,
    input  [15 : 0]     din32,
    input  [15 : 0]     din33,
    input  [15 : 0]     din34,
    input  [15 : 0]     din35,
    input  [15 : 0]     din36,
    input  [15 : 0]     din37,
    input  [15 : 0]     din38,
    input  [15 : 0]     din39,
    input  [15 : 0]     din40,
    input  [15 : 0]     din41,
    input  [15 : 0]     din42,
    input  [15 : 0]     din43,
    input  [15 : 0]     din44,
    input  [15 : 0]     din45,
    input  [15 : 0]     din46,
    input  [15 : 0]     din47,
    input  [15 : 0]     din48,
    input  [15 : 0]     din49,
    input  [15 : 0]     din50,
    input  [15 : 0]     din51,
    input  [15 : 0]     din52,
    input  [15 : 0]     din53,
    input  [15 : 0]     din54,
    input  [15 : 0]     din55,
    input  [15 : 0]     din56,
    input  [15 : 0]     din57,
    input  [15 : 0]     din58,
    input  [15 : 0]     din59,
    input  [15 : 0]     din60,
    input  [15 : 0]     din61,
    input  [15 : 0]     din62,
    input  [15 : 0]     din63,
    input  [15 : 0]     din64,
    input  [15 : 0]     din65,
    input  [15 : 0]     din66,
    input  [15 : 0]     din67,
    input  [15 : 0]     din68,
    input  [15 : 0]     din69,
    input  [15 : 0]     din70,
    input  [15 : 0]     din71,
    input  [15 : 0]     din72,
    input  [15 : 0]     din73,
    input  [15 : 0]     din74,
    input  [15 : 0]     din75,
    input  [15 : 0]     din76,
    input  [15 : 0]     din77,
    input  [15 : 0]     din78,
    input  [15 : 0]     din79,
    input  [15 : 0]     din80,
    input  [15 : 0]     din81,
    input  [15 : 0]     din82,
    input  [15 : 0]     din83,
    input  [15 : 0]     din84,
    input  [15 : 0]     din85,
    input  [15 : 0]     din86,
    input  [15 : 0]     din87,
    input  [15 : 0]     din88,
    input  [15 : 0]     din89,
    input  [15 : 0]     din90,
    input  [15 : 0]     din91,
    input  [15 : 0]     din92,
    input  [15 : 0]     din93,
    input  [15 : 0]     din94,
    input  [15 : 0]     din95,
    input  [15 : 0]     din96,
    input  [15 : 0]     din97,
    input  [15 : 0]     din98,
    input  [15 : 0]     din99,
    input  [15 : 0]     din100,
    input  [15 : 0]     din101,
    input  [15 : 0]     din102,
    input  [15 : 0]     din103,
    input  [15 : 0]     din104,
    input  [15 : 0]     din105,
    input  [15 : 0]     din106,
    input  [15 : 0]     din107,
    input  [15 : 0]     din108,
    input  [15 : 0]     din109,
    input  [15 : 0]     din110,
    input  [15 : 0]     din111,
    input  [15 : 0]     din112,
    input  [15 : 0]     din113,
    input  [15 : 0]     din114,
    input  [15 : 0]     din115,
    input  [15 : 0]     din116,
    input  [15 : 0]     din117,
    input  [15 : 0]     din118,
    input  [15 : 0]     din119,
    input  [15 : 0]     din120,
    input  [15 : 0]     din121,
    input  [15 : 0]     din122,
    input  [15 : 0]     din123,
    input  [15 : 0]     din124,
    input  [15 : 0]     din125,
    input  [15 : 0]     din126,
    input  [15 : 0]     din127,
    input  [15 : 0]     din128,
    input  [15 : 0]     din129,
    input  [15 : 0]     din130,
    input  [15 : 0]     din131,
    input  [15 : 0]     din132,
    input  [15 : 0]     din133,
    input  [15 : 0]     din134,
    input  [15 : 0]     din135,
    input  [15 : 0]     din136,
    input  [15 : 0]     din137,
    input  [15 : 0]     din138,
    input  [15 : 0]     din139,
    input  [15 : 0]     din140,
    input  [15 : 0]     din141,
    input  [15 : 0]     din142,
    input  [15 : 0]     din143,
    input  [15 : 0]     din144,
    input  [15 : 0]     din145,
    input  [15 : 0]     din146,
    input  [15 : 0]     din147,
    input  [15 : 0]     din148,
    input  [15 : 0]     din149,
    input  [15 : 0]     din150,
    input  [15 : 0]     din151,
    input  [15 : 0]     din152,
    input  [15 : 0]     din153,
    input  [15 : 0]     din154,
    input  [15 : 0]     din155,
    input  [15 : 0]     din156,
    input  [15 : 0]     din157,
    input  [15 : 0]     din158,
    input  [15 : 0]     din159,
    input  [15 : 0]     din160,
    input  [15 : 0]     din161,
    input  [15 : 0]     din162,
    input  [15 : 0]     din163,
    input  [15 : 0]     din164,
    input  [15 : 0]     din165,
    input  [15 : 0]     din166,
    input  [15 : 0]     din167,
    input  [15 : 0]     din168,
    input  [15 : 0]     din169,
    input  [15 : 0]     din170,
    input  [15 : 0]     din171,
    input  [15 : 0]     din172,
    input  [15 : 0]     din173,
    input  [15 : 0]     din174,
    input  [15 : 0]     din175,
    input  [15 : 0]     din176,
    input  [15 : 0]     din177,
    input  [15 : 0]     din178,
    input  [15 : 0]     din179,
    input  [15 : 0]     din180,
    input  [15 : 0]     din181,
    input  [15 : 0]     din182,
    input  [15 : 0]     din183,
    input  [15 : 0]     din184,
    input  [15 : 0]     din185,
    input  [15 : 0]     din186,
    input  [15 : 0]     din187,
    input  [15 : 0]     din188,
    input  [15 : 0]     din189,
    input  [15 : 0]     din190,
    input  [15 : 0]     din191,
    input  [15 : 0]     din192,
    input  [15 : 0]     din193,
    input  [15 : 0]     din194,
    input  [15 : 0]     din195,
    input  [15 : 0]     din196,
    input  [15 : 0]     din197,
    input  [15 : 0]     din198,
    input  [15 : 0]     din199,
    input  [15 : 0]     din200,
    input  [15 : 0]     din201,
    input  [15 : 0]     din202,
    input  [15 : 0]     din203,
    input  [15 : 0]     din204,
    input  [15 : 0]     din205,
    input  [15 : 0]     din206,
    input  [15 : 0]     din207,
    input  [15 : 0]     din208,
    input  [15 : 0]     din209,
    input  [15 : 0]     din210,
    input  [15 : 0]     din211,
    input  [15 : 0]     din212,
    input  [15 : 0]     din213,
    input  [15 : 0]     din214,
    input  [15 : 0]     din215,
    input  [15 : 0]     din216,
    input  [15 : 0]     din217,
    input  [15 : 0]     din218,
    input  [15 : 0]     din219,
    input  [15 : 0]     din220,
    input  [15 : 0]     din221,
    input  [15 : 0]     din222,
    input  [15 : 0]     din223,
    input  [15 : 0]     din224,
    input  [15 : 0]     din225,
    input  [15 : 0]     din226,
    input  [15 : 0]     din227,
    input  [15 : 0]     din228,
    input  [15 : 0]     din229,
    input  [15 : 0]     din230,
    input  [15 : 0]     din231,
    input  [15 : 0]     din232,
    input  [15 : 0]     din233,
    input  [15 : 0]     din234,
    input  [15 : 0]     din235,
    input  [15 : 0]     din236,
    input  [15 : 0]     din237,
    input  [15 : 0]     din238,
    input  [15 : 0]     din239,
    input  [15 : 0]     din240,
    input  [15 : 0]     din241,
    input  [15 : 0]     din242,
    input  [15 : 0]     din243,
    input  [15 : 0]     din244,
    input  [15 : 0]     din245,
    input  [15 : 0]     din246,
    input  [15 : 0]     din247,
    input  [15 : 0]     din248,
    input  [15 : 0]     din249,
    input  [15 : 0]     din250,
    input  [15 : 0]     din251,
    input  [15 : 0]     din252,
    input  [15 : 0]     din253,
    input  [15 : 0]     din254,
    input  [15 : 0]     din255,
    input  [15 : 0]     din256,
    input  [15 : 0]     din257,
    input  [15 : 0]     din258,
    input  [15 : 0]     din259,
    input  [15 : 0]     din260,
    input  [15 : 0]     din261,
    input  [15 : 0]     din262,
    input  [15 : 0]     din263,
    input  [15 : 0]     din264,
    input  [15 : 0]     din265,
    input  [15 : 0]     din266,
    input  [15 : 0]     din267,
    input  [15 : 0]     din268,
    input  [15 : 0]     din269,
    input  [15 : 0]     din270,
    input  [15 : 0]     din271,
    input  [15 : 0]     din272,
    input  [15 : 0]     din273,
    input  [15 : 0]     din274,
    input  [15 : 0]     din275,
    input  [15 : 0]     din276,
    input  [15 : 0]     din277,
    input  [15 : 0]     din278,
    input  [15 : 0]     din279,
    input  [15 : 0]     din280,
    input  [15 : 0]     din281,
    input  [15 : 0]     din282,
    input  [15 : 0]     din283,
    input  [15 : 0]     din284,
    input  [15 : 0]     din285,
    input  [15 : 0]     din286,
    input  [15 : 0]     din287,
    input  [15 : 0]     din288,
    input  [15 : 0]     din289,
    input  [15 : 0]     din290,
    input  [15 : 0]     din291,
    input  [15 : 0]     din292,
    input  [15 : 0]     din293,
    input  [15 : 0]     din294,
    input  [15 : 0]     din295,
    input  [15 : 0]     din296,
    input  [15 : 0]     din297,
    input  [15 : 0]     din298,
    input  [15 : 0]     din299,
    input  [15 : 0]     din300,
    input  [15 : 0]     din301,
    input  [15 : 0]     din302,
    input  [15 : 0]     din303,
    input  [15 : 0]     din304,
    input  [15 : 0]     din305,
    input  [15 : 0]     din306,
    input  [15 : 0]     din307,
    input  [15 : 0]     din308,
    input  [15 : 0]     din309,
    input  [15 : 0]     din310,
    input  [15 : 0]     din311,
    input  [15 : 0]     din312,
    input  [15 : 0]     din313,
    input  [15 : 0]     din314,
    input  [15 : 0]     din315,
    input  [15 : 0]     din316,
    input  [15 : 0]     din317,
    input  [15 : 0]     din318,
    input  [15 : 0]     din319,
    input  [15 : 0]     din320,
    input  [15 : 0]     din321,
    input  [15 : 0]     din322,
    input  [15 : 0]     din323,
    input  [15 : 0]     din324,
    input  [15 : 0]     din325,
    input  [15 : 0]     din326,
    input  [15 : 0]     din327,
    input  [15 : 0]     din328,
    input  [15 : 0]     din329,
    input  [15 : 0]     din330,
    input  [15 : 0]     din331,
    input  [15 : 0]     din332,
    input  [15 : 0]     din333,
    input  [15 : 0]     din334,
    input  [15 : 0]     din335,
    input  [15 : 0]     din336,
    input  [15 : 0]     din337,
    input  [15 : 0]     din338,
    input  [15 : 0]     din339,
    input  [15 : 0]     din340,
    input  [15 : 0]     din341,
    input  [15 : 0]     din342,
    input  [15 : 0]     din343,
    input  [15 : 0]     din344,
    input  [15 : 0]     din345,
    input  [15 : 0]     din346,
    input  [15 : 0]     din347,
    input  [15 : 0]     din348,
    input  [15 : 0]     din349,
    input  [15 : 0]     din350,
    input  [15 : 0]     din351,
    input  [15 : 0]     din352,
    input  [15 : 0]     din353,
    input  [15 : 0]     din354,
    input  [15 : 0]     din355,
    input  [15 : 0]     din356,
    input  [15 : 0]     din357,
    input  [15 : 0]     din358,
    input  [15 : 0]     din359,
    input  [15 : 0]     din360,
    input  [15 : 0]     din361,
    input  [15 : 0]     din362,
    input  [15 : 0]     din363,
    input  [15 : 0]     din364,
    input  [15 : 0]     din365,
    input  [15 : 0]     din366,
    input  [15 : 0]     din367,
    input  [15 : 0]     din368,
    input  [15 : 0]     din369,
    input  [15 : 0]     din370,
    input  [15 : 0]     din371,
    input  [15 : 0]     din372,
    input  [15 : 0]     din373,
    input  [15 : 0]     din374,
    input  [15 : 0]     din375,
    input  [15 : 0]     din376,
    input  [15 : 0]     din377,
    input  [15 : 0]     din378,
    input  [15 : 0]     din379,
    input  [15 : 0]     din380,
    input  [15 : 0]     din381,
    input  [15 : 0]     din382,
    input  [15 : 0]     din383,
    input  [15 : 0]     din384,
    input  [15 : 0]     din385,
    input  [15 : 0]     din386,
    input  [15 : 0]     din387,
    input  [15 : 0]     din388,
    input  [15 : 0]     din389,
    input  [15 : 0]     din390,
    input  [15 : 0]     din391,
    input  [15 : 0]     din392,
    input  [15 : 0]     din393,
    input  [15 : 0]     din394,
    input  [15 : 0]     din395,
    input  [15 : 0]     din396,
    input  [15 : 0]     din397,
    input  [15 : 0]     din398,
    input  [15 : 0]     din399,
    input  [15 : 0]     din400,
    input  [15 : 0]     din401,
    input  [15 : 0]     din402,
    input  [15 : 0]     din403,
    input  [15 : 0]     din404,
    input  [15 : 0]     din405,
    input  [15 : 0]     din406,
    input  [15 : 0]     din407,
    input  [15 : 0]     din408,
    input  [15 : 0]     din409,
    input  [15 : 0]     din410,
    input  [15 : 0]     din411,
    input  [15 : 0]     din412,
    input  [15 : 0]     din413,
    input  [15 : 0]     din414,
    input  [15 : 0]     din415,
    input  [15 : 0]     din416,
    input  [15 : 0]     din417,
    input  [15 : 0]     din418,
    input  [15 : 0]     din419,
    input  [15 : 0]     din420,
    input  [15 : 0]     din421,
    input  [15 : 0]     din422,
    input  [15 : 0]     din423,
    input  [15 : 0]     din424,
    input  [15 : 0]     din425,
    input  [15 : 0]     din426,
    input  [15 : 0]     din427,
    input  [15 : 0]     din428,
    input  [15 : 0]     din429,
    input  [15 : 0]     din430,
    input  [15 : 0]     din431,
    input  [15 : 0]     din432,
    input  [15 : 0]     din433,
    input  [15 : 0]     din434,
    input  [15 : 0]     din435,
    input  [15 : 0]     din436,
    input  [15 : 0]     din437,
    input  [15 : 0]     din438,
    input  [15 : 0]     din439,
    input  [15 : 0]     din440,
    input  [15 : 0]     din441,
    input  [15 : 0]     din442,
    input  [15 : 0]     din443,
    input  [15 : 0]     din444,
    input  [15 : 0]     din445,
    input  [15 : 0]     din446,
    input  [15 : 0]     din447,
    input  [15 : 0]     din448,
    input  [15 : 0]     din449,
    input  [15 : 0]     din450,
    input  [15 : 0]     din451,
    input  [15 : 0]     din452,
    input  [15 : 0]     din453,
    input  [15 : 0]     din454,
    input  [15 : 0]     din455,
    input  [15 : 0]     din456,
    input  [15 : 0]     din457,
    input  [15 : 0]     din458,
    input  [15 : 0]     din459,
    input  [15 : 0]     din460,
    input  [15 : 0]     din461,
    input  [15 : 0]     din462,
    input  [15 : 0]     din463,
    input  [15 : 0]     din464,
    input  [15 : 0]     din465,
    input  [15 : 0]     din466,
    input  [15 : 0]     din467,
    input  [15 : 0]     din468,
    input  [15 : 0]     din469,
    input  [15 : 0]     din470,
    input  [15 : 0]     din471,
    input  [15 : 0]     din472,
    input  [15 : 0]     din473,
    input  [15 : 0]     din474,
    input  [15 : 0]     din475,
    input  [15 : 0]     din476,
    input  [15 : 0]     din477,
    input  [15 : 0]     din478,
    input  [15 : 0]     din479,
    input  [15 : 0]     din480,
    input  [15 : 0]     din481,
    input  [15 : 0]     din482,
    input  [15 : 0]     din483,
    input  [15 : 0]     din484,
    input  [15 : 0]     din485,
    input  [15 : 0]     din486,
    input  [15 : 0]     din487,
    input  [15 : 0]     din488,
    input  [15 : 0]     din489,
    input  [15 : 0]     din490,
    input  [15 : 0]     din491,
    input  [15 : 0]     din492,
    input  [15 : 0]     din493,
    input  [15 : 0]     din494,
    input  [15 : 0]     din495,
    input  [15 : 0]     din496,
    input  [15 : 0]     din497,
    input  [15 : 0]     din498,
    input  [15 : 0]     din499,
    input  [15 : 0]     din500,
    input  [15 : 0]     din501,
    input  [15 : 0]     din502,
    input  [15 : 0]     din503,
    input  [15 : 0]     din504,
    input  [15 : 0]     din505,
    input  [15 : 0]     din506,
    input  [15 : 0]     din507,
    input  [15 : 0]     din508,
    input  [15 : 0]     din509,
    input  [15 : 0]     din510,
    input  [15 : 0]     din511,
    input  [15 : 0]     din512,
    input  [15 : 0]     din513,
    input  [15 : 0]     din514,
    input  [15 : 0]     din515,
    input  [15 : 0]     din516,
    input  [15 : 0]     din517,
    input  [15 : 0]     din518,
    input  [15 : 0]     din519,
    input  [15 : 0]     din520,
    input  [15 : 0]     din521,
    input  [15 : 0]     din522,
    input  [15 : 0]     din523,
    input  [15 : 0]     din524,
    input  [15 : 0]     din525,
    input  [15 : 0]     din526,
    input  [15 : 0]     din527,
    input  [15 : 0]     din528,
    input  [15 : 0]     din529,
    input  [15 : 0]     din530,
    input  [15 : 0]     din531,
    input  [15 : 0]     din532,
    input  [15 : 0]     din533,
    input  [15 : 0]     din534,
    input  [15 : 0]     din535,
    input  [15 : 0]     din536,
    input  [15 : 0]     din537,
    input  [15 : 0]     din538,
    input  [15 : 0]     din539,
    input  [15 : 0]     din540,
    input  [15 : 0]     din541,
    input  [15 : 0]     din542,
    input  [15 : 0]     din543,
    input  [15 : 0]     din544,
    input  [15 : 0]     din545,
    input  [15 : 0]     din546,
    input  [15 : 0]     din547,
    input  [15 : 0]     din548,
    input  [15 : 0]     din549,
    input  [15 : 0]     din550,
    input  [15 : 0]     din551,
    input  [15 : 0]     din552,
    input  [15 : 0]     din553,
    input  [15 : 0]     din554,
    input  [15 : 0]     din555,
    input  [15 : 0]     din556,
    input  [15 : 0]     din557,
    input  [15 : 0]     din558,
    input  [15 : 0]     din559,
    input  [15 : 0]     din560,
    input  [15 : 0]     din561,
    input  [15 : 0]     din562,
    input  [15 : 0]     din563,
    input  [15 : 0]     din564,
    input  [15 : 0]     din565,
    input  [15 : 0]     din566,
    input  [15 : 0]     din567,
    input  [15 : 0]     din568,
    input  [15 : 0]     din569,
    input  [15 : 0]     din570,
    input  [15 : 0]     din571,
    input  [15 : 0]     din572,
    input  [15 : 0]     din573,
    input  [15 : 0]     din574,
    input  [15 : 0]     din575,
    input  [9 : 0]    din576,
    output [15 : 0]   dout);

// puts internal signals
wire [9 : 0]     sel;
// level 1 signals
wire [15 : 0]         mux_1_0;
wire [15 : 0]         mux_1_1;
wire [15 : 0]         mux_1_2;
wire [15 : 0]         mux_1_3;
wire [15 : 0]         mux_1_4;
wire [15 : 0]         mux_1_5;
wire [15 : 0]         mux_1_6;
wire [15 : 0]         mux_1_7;
wire [15 : 0]         mux_1_8;
wire [15 : 0]         mux_1_9;
wire [15 : 0]         mux_1_10;
wire [15 : 0]         mux_1_11;
wire [15 : 0]         mux_1_12;
wire [15 : 0]         mux_1_13;
wire [15 : 0]         mux_1_14;
wire [15 : 0]         mux_1_15;
wire [15 : 0]         mux_1_16;
wire [15 : 0]         mux_1_17;
wire [15 : 0]         mux_1_18;
wire [15 : 0]         mux_1_19;
wire [15 : 0]         mux_1_20;
wire [15 : 0]         mux_1_21;
wire [15 : 0]         mux_1_22;
wire [15 : 0]         mux_1_23;
wire [15 : 0]         mux_1_24;
wire [15 : 0]         mux_1_25;
wire [15 : 0]         mux_1_26;
wire [15 : 0]         mux_1_27;
wire [15 : 0]         mux_1_28;
wire [15 : 0]         mux_1_29;
wire [15 : 0]         mux_1_30;
wire [15 : 0]         mux_1_31;
wire [15 : 0]         mux_1_32;
wire [15 : 0]         mux_1_33;
wire [15 : 0]         mux_1_34;
wire [15 : 0]         mux_1_35;
wire [15 : 0]         mux_1_36;
wire [15 : 0]         mux_1_37;
wire [15 : 0]         mux_1_38;
wire [15 : 0]         mux_1_39;
wire [15 : 0]         mux_1_40;
wire [15 : 0]         mux_1_41;
wire [15 : 0]         mux_1_42;
wire [15 : 0]         mux_1_43;
wire [15 : 0]         mux_1_44;
wire [15 : 0]         mux_1_45;
wire [15 : 0]         mux_1_46;
wire [15 : 0]         mux_1_47;
wire [15 : 0]         mux_1_48;
wire [15 : 0]         mux_1_49;
wire [15 : 0]         mux_1_50;
wire [15 : 0]         mux_1_51;
wire [15 : 0]         mux_1_52;
wire [15 : 0]         mux_1_53;
wire [15 : 0]         mux_1_54;
wire [15 : 0]         mux_1_55;
wire [15 : 0]         mux_1_56;
wire [15 : 0]         mux_1_57;
wire [15 : 0]         mux_1_58;
wire [15 : 0]         mux_1_59;
wire [15 : 0]         mux_1_60;
wire [15 : 0]         mux_1_61;
wire [15 : 0]         mux_1_62;
wire [15 : 0]         mux_1_63;
wire [15 : 0]         mux_1_64;
wire [15 : 0]         mux_1_65;
wire [15 : 0]         mux_1_66;
wire [15 : 0]         mux_1_67;
wire [15 : 0]         mux_1_68;
wire [15 : 0]         mux_1_69;
wire [15 : 0]         mux_1_70;
wire [15 : 0]         mux_1_71;
wire [15 : 0]         mux_1_72;
wire [15 : 0]         mux_1_73;
wire [15 : 0]         mux_1_74;
wire [15 : 0]         mux_1_75;
wire [15 : 0]         mux_1_76;
wire [15 : 0]         mux_1_77;
wire [15 : 0]         mux_1_78;
wire [15 : 0]         mux_1_79;
wire [15 : 0]         mux_1_80;
wire [15 : 0]         mux_1_81;
wire [15 : 0]         mux_1_82;
wire [15 : 0]         mux_1_83;
wire [15 : 0]         mux_1_84;
wire [15 : 0]         mux_1_85;
wire [15 : 0]         mux_1_86;
wire [15 : 0]         mux_1_87;
wire [15 : 0]         mux_1_88;
wire [15 : 0]         mux_1_89;
wire [15 : 0]         mux_1_90;
wire [15 : 0]         mux_1_91;
wire [15 : 0]         mux_1_92;
wire [15 : 0]         mux_1_93;
wire [15 : 0]         mux_1_94;
wire [15 : 0]         mux_1_95;
wire [15 : 0]         mux_1_96;
wire [15 : 0]         mux_1_97;
wire [15 : 0]         mux_1_98;
wire [15 : 0]         mux_1_99;
wire [15 : 0]         mux_1_100;
wire [15 : 0]         mux_1_101;
wire [15 : 0]         mux_1_102;
wire [15 : 0]         mux_1_103;
wire [15 : 0]         mux_1_104;
wire [15 : 0]         mux_1_105;
wire [15 : 0]         mux_1_106;
wire [15 : 0]         mux_1_107;
wire [15 : 0]         mux_1_108;
wire [15 : 0]         mux_1_109;
wire [15 : 0]         mux_1_110;
wire [15 : 0]         mux_1_111;
wire [15 : 0]         mux_1_112;
wire [15 : 0]         mux_1_113;
wire [15 : 0]         mux_1_114;
wire [15 : 0]         mux_1_115;
wire [15 : 0]         mux_1_116;
wire [15 : 0]         mux_1_117;
wire [15 : 0]         mux_1_118;
wire [15 : 0]         mux_1_119;
wire [15 : 0]         mux_1_120;
wire [15 : 0]         mux_1_121;
wire [15 : 0]         mux_1_122;
wire [15 : 0]         mux_1_123;
wire [15 : 0]         mux_1_124;
wire [15 : 0]         mux_1_125;
wire [15 : 0]         mux_1_126;
wire [15 : 0]         mux_1_127;
wire [15 : 0]         mux_1_128;
wire [15 : 0]         mux_1_129;
wire [15 : 0]         mux_1_130;
wire [15 : 0]         mux_1_131;
wire [15 : 0]         mux_1_132;
wire [15 : 0]         mux_1_133;
wire [15 : 0]         mux_1_134;
wire [15 : 0]         mux_1_135;
wire [15 : 0]         mux_1_136;
wire [15 : 0]         mux_1_137;
wire [15 : 0]         mux_1_138;
wire [15 : 0]         mux_1_139;
wire [15 : 0]         mux_1_140;
wire [15 : 0]         mux_1_141;
wire [15 : 0]         mux_1_142;
wire [15 : 0]         mux_1_143;
wire [15 : 0]         mux_1_144;
wire [15 : 0]         mux_1_145;
wire [15 : 0]         mux_1_146;
wire [15 : 0]         mux_1_147;
wire [15 : 0]         mux_1_148;
wire [15 : 0]         mux_1_149;
wire [15 : 0]         mux_1_150;
wire [15 : 0]         mux_1_151;
wire [15 : 0]         mux_1_152;
wire [15 : 0]         mux_1_153;
wire [15 : 0]         mux_1_154;
wire [15 : 0]         mux_1_155;
wire [15 : 0]         mux_1_156;
wire [15 : 0]         mux_1_157;
wire [15 : 0]         mux_1_158;
wire [15 : 0]         mux_1_159;
wire [15 : 0]         mux_1_160;
wire [15 : 0]         mux_1_161;
wire [15 : 0]         mux_1_162;
wire [15 : 0]         mux_1_163;
wire [15 : 0]         mux_1_164;
wire [15 : 0]         mux_1_165;
wire [15 : 0]         mux_1_166;
wire [15 : 0]         mux_1_167;
wire [15 : 0]         mux_1_168;
wire [15 : 0]         mux_1_169;
wire [15 : 0]         mux_1_170;
wire [15 : 0]         mux_1_171;
wire [15 : 0]         mux_1_172;
wire [15 : 0]         mux_1_173;
wire [15 : 0]         mux_1_174;
wire [15 : 0]         mux_1_175;
wire [15 : 0]         mux_1_176;
wire [15 : 0]         mux_1_177;
wire [15 : 0]         mux_1_178;
wire [15 : 0]         mux_1_179;
wire [15 : 0]         mux_1_180;
wire [15 : 0]         mux_1_181;
wire [15 : 0]         mux_1_182;
wire [15 : 0]         mux_1_183;
wire [15 : 0]         mux_1_184;
wire [15 : 0]         mux_1_185;
wire [15 : 0]         mux_1_186;
wire [15 : 0]         mux_1_187;
wire [15 : 0]         mux_1_188;
wire [15 : 0]         mux_1_189;
wire [15 : 0]         mux_1_190;
wire [15 : 0]         mux_1_191;
wire [15 : 0]         mux_1_192;
wire [15 : 0]         mux_1_193;
wire [15 : 0]         mux_1_194;
wire [15 : 0]         mux_1_195;
wire [15 : 0]         mux_1_196;
wire [15 : 0]         mux_1_197;
wire [15 : 0]         mux_1_198;
wire [15 : 0]         mux_1_199;
wire [15 : 0]         mux_1_200;
wire [15 : 0]         mux_1_201;
wire [15 : 0]         mux_1_202;
wire [15 : 0]         mux_1_203;
wire [15 : 0]         mux_1_204;
wire [15 : 0]         mux_1_205;
wire [15 : 0]         mux_1_206;
wire [15 : 0]         mux_1_207;
wire [15 : 0]         mux_1_208;
wire [15 : 0]         mux_1_209;
wire [15 : 0]         mux_1_210;
wire [15 : 0]         mux_1_211;
wire [15 : 0]         mux_1_212;
wire [15 : 0]         mux_1_213;
wire [15 : 0]         mux_1_214;
wire [15 : 0]         mux_1_215;
wire [15 : 0]         mux_1_216;
wire [15 : 0]         mux_1_217;
wire [15 : 0]         mux_1_218;
wire [15 : 0]         mux_1_219;
wire [15 : 0]         mux_1_220;
wire [15 : 0]         mux_1_221;
wire [15 : 0]         mux_1_222;
wire [15 : 0]         mux_1_223;
wire [15 : 0]         mux_1_224;
wire [15 : 0]         mux_1_225;
wire [15 : 0]         mux_1_226;
wire [15 : 0]         mux_1_227;
wire [15 : 0]         mux_1_228;
wire [15 : 0]         mux_1_229;
wire [15 : 0]         mux_1_230;
wire [15 : 0]         mux_1_231;
wire [15 : 0]         mux_1_232;
wire [15 : 0]         mux_1_233;
wire [15 : 0]         mux_1_234;
wire [15 : 0]         mux_1_235;
wire [15 : 0]         mux_1_236;
wire [15 : 0]         mux_1_237;
wire [15 : 0]         mux_1_238;
wire [15 : 0]         mux_1_239;
wire [15 : 0]         mux_1_240;
wire [15 : 0]         mux_1_241;
wire [15 : 0]         mux_1_242;
wire [15 : 0]         mux_1_243;
wire [15 : 0]         mux_1_244;
wire [15 : 0]         mux_1_245;
wire [15 : 0]         mux_1_246;
wire [15 : 0]         mux_1_247;
wire [15 : 0]         mux_1_248;
wire [15 : 0]         mux_1_249;
wire [15 : 0]         mux_1_250;
wire [15 : 0]         mux_1_251;
wire [15 : 0]         mux_1_252;
wire [15 : 0]         mux_1_253;
wire [15 : 0]         mux_1_254;
wire [15 : 0]         mux_1_255;
wire [15 : 0]         mux_1_256;
wire [15 : 0]         mux_1_257;
wire [15 : 0]         mux_1_258;
wire [15 : 0]         mux_1_259;
wire [15 : 0]         mux_1_260;
wire [15 : 0]         mux_1_261;
wire [15 : 0]         mux_1_262;
wire [15 : 0]         mux_1_263;
wire [15 : 0]         mux_1_264;
wire [15 : 0]         mux_1_265;
wire [15 : 0]         mux_1_266;
wire [15 : 0]         mux_1_267;
wire [15 : 0]         mux_1_268;
wire [15 : 0]         mux_1_269;
wire [15 : 0]         mux_1_270;
wire [15 : 0]         mux_1_271;
wire [15 : 0]         mux_1_272;
wire [15 : 0]         mux_1_273;
wire [15 : 0]         mux_1_274;
wire [15 : 0]         mux_1_275;
wire [15 : 0]         mux_1_276;
wire [15 : 0]         mux_1_277;
wire [15 : 0]         mux_1_278;
wire [15 : 0]         mux_1_279;
wire [15 : 0]         mux_1_280;
wire [15 : 0]         mux_1_281;
wire [15 : 0]         mux_1_282;
wire [15 : 0]         mux_1_283;
wire [15 : 0]         mux_1_284;
wire [15 : 0]         mux_1_285;
wire [15 : 0]         mux_1_286;
wire [15 : 0]         mux_1_287;
// level 2 signals
wire [15 : 0]         mux_2_0;
wire [15 : 0]         mux_2_1;
wire [15 : 0]         mux_2_2;
wire [15 : 0]         mux_2_3;
wire [15 : 0]         mux_2_4;
wire [15 : 0]         mux_2_5;
wire [15 : 0]         mux_2_6;
wire [15 : 0]         mux_2_7;
wire [15 : 0]         mux_2_8;
wire [15 : 0]         mux_2_9;
wire [15 : 0]         mux_2_10;
wire [15 : 0]         mux_2_11;
wire [15 : 0]         mux_2_12;
wire [15 : 0]         mux_2_13;
wire [15 : 0]         mux_2_14;
wire [15 : 0]         mux_2_15;
wire [15 : 0]         mux_2_16;
wire [15 : 0]         mux_2_17;
wire [15 : 0]         mux_2_18;
wire [15 : 0]         mux_2_19;
wire [15 : 0]         mux_2_20;
wire [15 : 0]         mux_2_21;
wire [15 : 0]         mux_2_22;
wire [15 : 0]         mux_2_23;
wire [15 : 0]         mux_2_24;
wire [15 : 0]         mux_2_25;
wire [15 : 0]         mux_2_26;
wire [15 : 0]         mux_2_27;
wire [15 : 0]         mux_2_28;
wire [15 : 0]         mux_2_29;
wire [15 : 0]         mux_2_30;
wire [15 : 0]         mux_2_31;
wire [15 : 0]         mux_2_32;
wire [15 : 0]         mux_2_33;
wire [15 : 0]         mux_2_34;
wire [15 : 0]         mux_2_35;
wire [15 : 0]         mux_2_36;
wire [15 : 0]         mux_2_37;
wire [15 : 0]         mux_2_38;
wire [15 : 0]         mux_2_39;
wire [15 : 0]         mux_2_40;
wire [15 : 0]         mux_2_41;
wire [15 : 0]         mux_2_42;
wire [15 : 0]         mux_2_43;
wire [15 : 0]         mux_2_44;
wire [15 : 0]         mux_2_45;
wire [15 : 0]         mux_2_46;
wire [15 : 0]         mux_2_47;
wire [15 : 0]         mux_2_48;
wire [15 : 0]         mux_2_49;
wire [15 : 0]         mux_2_50;
wire [15 : 0]         mux_2_51;
wire [15 : 0]         mux_2_52;
wire [15 : 0]         mux_2_53;
wire [15 : 0]         mux_2_54;
wire [15 : 0]         mux_2_55;
wire [15 : 0]         mux_2_56;
wire [15 : 0]         mux_2_57;
wire [15 : 0]         mux_2_58;
wire [15 : 0]         mux_2_59;
wire [15 : 0]         mux_2_60;
wire [15 : 0]         mux_2_61;
wire [15 : 0]         mux_2_62;
wire [15 : 0]         mux_2_63;
wire [15 : 0]         mux_2_64;
wire [15 : 0]         mux_2_65;
wire [15 : 0]         mux_2_66;
wire [15 : 0]         mux_2_67;
wire [15 : 0]         mux_2_68;
wire [15 : 0]         mux_2_69;
wire [15 : 0]         mux_2_70;
wire [15 : 0]         mux_2_71;
wire [15 : 0]         mux_2_72;
wire [15 : 0]         mux_2_73;
wire [15 : 0]         mux_2_74;
wire [15 : 0]         mux_2_75;
wire [15 : 0]         mux_2_76;
wire [15 : 0]         mux_2_77;
wire [15 : 0]         mux_2_78;
wire [15 : 0]         mux_2_79;
wire [15 : 0]         mux_2_80;
wire [15 : 0]         mux_2_81;
wire [15 : 0]         mux_2_82;
wire [15 : 0]         mux_2_83;
wire [15 : 0]         mux_2_84;
wire [15 : 0]         mux_2_85;
wire [15 : 0]         mux_2_86;
wire [15 : 0]         mux_2_87;
wire [15 : 0]         mux_2_88;
wire [15 : 0]         mux_2_89;
wire [15 : 0]         mux_2_90;
wire [15 : 0]         mux_2_91;
wire [15 : 0]         mux_2_92;
wire [15 : 0]         mux_2_93;
wire [15 : 0]         mux_2_94;
wire [15 : 0]         mux_2_95;
wire [15 : 0]         mux_2_96;
wire [15 : 0]         mux_2_97;
wire [15 : 0]         mux_2_98;
wire [15 : 0]         mux_2_99;
wire [15 : 0]         mux_2_100;
wire [15 : 0]         mux_2_101;
wire [15 : 0]         mux_2_102;
wire [15 : 0]         mux_2_103;
wire [15 : 0]         mux_2_104;
wire [15 : 0]         mux_2_105;
wire [15 : 0]         mux_2_106;
wire [15 : 0]         mux_2_107;
wire [15 : 0]         mux_2_108;
wire [15 : 0]         mux_2_109;
wire [15 : 0]         mux_2_110;
wire [15 : 0]         mux_2_111;
wire [15 : 0]         mux_2_112;
wire [15 : 0]         mux_2_113;
wire [15 : 0]         mux_2_114;
wire [15 : 0]         mux_2_115;
wire [15 : 0]         mux_2_116;
wire [15 : 0]         mux_2_117;
wire [15 : 0]         mux_2_118;
wire [15 : 0]         mux_2_119;
wire [15 : 0]         mux_2_120;
wire [15 : 0]         mux_2_121;
wire [15 : 0]         mux_2_122;
wire [15 : 0]         mux_2_123;
wire [15 : 0]         mux_2_124;
wire [15 : 0]         mux_2_125;
wire [15 : 0]         mux_2_126;
wire [15 : 0]         mux_2_127;
wire [15 : 0]         mux_2_128;
wire [15 : 0]         mux_2_129;
wire [15 : 0]         mux_2_130;
wire [15 : 0]         mux_2_131;
wire [15 : 0]         mux_2_132;
wire [15 : 0]         mux_2_133;
wire [15 : 0]         mux_2_134;
wire [15 : 0]         mux_2_135;
wire [15 : 0]         mux_2_136;
wire [15 : 0]         mux_2_137;
wire [15 : 0]         mux_2_138;
wire [15 : 0]         mux_2_139;
wire [15 : 0]         mux_2_140;
wire [15 : 0]         mux_2_141;
wire [15 : 0]         mux_2_142;
wire [15 : 0]         mux_2_143;
// level 3 signals
wire [15 : 0]         mux_3_0;
wire [15 : 0]         mux_3_1;
wire [15 : 0]         mux_3_2;
wire [15 : 0]         mux_3_3;
wire [15 : 0]         mux_3_4;
wire [15 : 0]         mux_3_5;
wire [15 : 0]         mux_3_6;
wire [15 : 0]         mux_3_7;
wire [15 : 0]         mux_3_8;
wire [15 : 0]         mux_3_9;
wire [15 : 0]         mux_3_10;
wire [15 : 0]         mux_3_11;
wire [15 : 0]         mux_3_12;
wire [15 : 0]         mux_3_13;
wire [15 : 0]         mux_3_14;
wire [15 : 0]         mux_3_15;
wire [15 : 0]         mux_3_16;
wire [15 : 0]         mux_3_17;
wire [15 : 0]         mux_3_18;
wire [15 : 0]         mux_3_19;
wire [15 : 0]         mux_3_20;
wire [15 : 0]         mux_3_21;
wire [15 : 0]         mux_3_22;
wire [15 : 0]         mux_3_23;
wire [15 : 0]         mux_3_24;
wire [15 : 0]         mux_3_25;
wire [15 : 0]         mux_3_26;
wire [15 : 0]         mux_3_27;
wire [15 : 0]         mux_3_28;
wire [15 : 0]         mux_3_29;
wire [15 : 0]         mux_3_30;
wire [15 : 0]         mux_3_31;
wire [15 : 0]         mux_3_32;
wire [15 : 0]         mux_3_33;
wire [15 : 0]         mux_3_34;
wire [15 : 0]         mux_3_35;
wire [15 : 0]         mux_3_36;
wire [15 : 0]         mux_3_37;
wire [15 : 0]         mux_3_38;
wire [15 : 0]         mux_3_39;
wire [15 : 0]         mux_3_40;
wire [15 : 0]         mux_3_41;
wire [15 : 0]         mux_3_42;
wire [15 : 0]         mux_3_43;
wire [15 : 0]         mux_3_44;
wire [15 : 0]         mux_3_45;
wire [15 : 0]         mux_3_46;
wire [15 : 0]         mux_3_47;
wire [15 : 0]         mux_3_48;
wire [15 : 0]         mux_3_49;
wire [15 : 0]         mux_3_50;
wire [15 : 0]         mux_3_51;
wire [15 : 0]         mux_3_52;
wire [15 : 0]         mux_3_53;
wire [15 : 0]         mux_3_54;
wire [15 : 0]         mux_3_55;
wire [15 : 0]         mux_3_56;
wire [15 : 0]         mux_3_57;
wire [15 : 0]         mux_3_58;
wire [15 : 0]         mux_3_59;
wire [15 : 0]         mux_3_60;
wire [15 : 0]         mux_3_61;
wire [15 : 0]         mux_3_62;
wire [15 : 0]         mux_3_63;
wire [15 : 0]         mux_3_64;
wire [15 : 0]         mux_3_65;
wire [15 : 0]         mux_3_66;
wire [15 : 0]         mux_3_67;
wire [15 : 0]         mux_3_68;
wire [15 : 0]         mux_3_69;
wire [15 : 0]         mux_3_70;
wire [15 : 0]         mux_3_71;
// level 4 signals
wire [15 : 0]         mux_4_0;
wire [15 : 0]         mux_4_1;
wire [15 : 0]         mux_4_2;
wire [15 : 0]         mux_4_3;
wire [15 : 0]         mux_4_4;
wire [15 : 0]         mux_4_5;
wire [15 : 0]         mux_4_6;
wire [15 : 0]         mux_4_7;
wire [15 : 0]         mux_4_8;
wire [15 : 0]         mux_4_9;
wire [15 : 0]         mux_4_10;
wire [15 : 0]         mux_4_11;
wire [15 : 0]         mux_4_12;
wire [15 : 0]         mux_4_13;
wire [15 : 0]         mux_4_14;
wire [15 : 0]         mux_4_15;
wire [15 : 0]         mux_4_16;
wire [15 : 0]         mux_4_17;
wire [15 : 0]         mux_4_18;
wire [15 : 0]         mux_4_19;
wire [15 : 0]         mux_4_20;
wire [15 : 0]         mux_4_21;
wire [15 : 0]         mux_4_22;
wire [15 : 0]         mux_4_23;
wire [15 : 0]         mux_4_24;
wire [15 : 0]         mux_4_25;
wire [15 : 0]         mux_4_26;
wire [15 : 0]         mux_4_27;
wire [15 : 0]         mux_4_28;
wire [15 : 0]         mux_4_29;
wire [15 : 0]         mux_4_30;
wire [15 : 0]         mux_4_31;
wire [15 : 0]         mux_4_32;
wire [15 : 0]         mux_4_33;
wire [15 : 0]         mux_4_34;
wire [15 : 0]         mux_4_35;
// level 5 signals
wire [15 : 0]         mux_5_0;
wire [15 : 0]         mux_5_1;
wire [15 : 0]         mux_5_2;
wire [15 : 0]         mux_5_3;
wire [15 : 0]         mux_5_4;
wire [15 : 0]         mux_5_5;
wire [15 : 0]         mux_5_6;
wire [15 : 0]         mux_5_7;
wire [15 : 0]         mux_5_8;
wire [15 : 0]         mux_5_9;
wire [15 : 0]         mux_5_10;
wire [15 : 0]         mux_5_11;
wire [15 : 0]         mux_5_12;
wire [15 : 0]         mux_5_13;
wire [15 : 0]         mux_5_14;
wire [15 : 0]         mux_5_15;
wire [15 : 0]         mux_5_16;
wire [15 : 0]         mux_5_17;
// level 6 signals
wire [15 : 0]         mux_6_0;
wire [15 : 0]         mux_6_1;
wire [15 : 0]         mux_6_2;
wire [15 : 0]         mux_6_3;
wire [15 : 0]         mux_6_4;
wire [15 : 0]         mux_6_5;
wire [15 : 0]         mux_6_6;
wire [15 : 0]         mux_6_7;
wire [15 : 0]         mux_6_8;
// level 7 signals
wire [15 : 0]         mux_7_0;
wire [15 : 0]         mux_7_1;
wire [15 : 0]         mux_7_2;
wire [15 : 0]         mux_7_3;
wire [15 : 0]         mux_7_4;
// level 8 signals
wire [15 : 0]         mux_8_0;
wire [15 : 0]         mux_8_1;
wire [15 : 0]         mux_8_2;
// level 9 signals
wire [15 : 0]         mux_9_0;
wire [15 : 0]         mux_9_1;
// level 10 signals
wire [15 : 0]         mux_10_0;

assign sel = din576;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;
assign mux_1_2 = (sel[0] == 0)? din4 : din5;
assign mux_1_3 = (sel[0] == 0)? din6 : din7;
assign mux_1_4 = (sel[0] == 0)? din8 : din9;
assign mux_1_5 = (sel[0] == 0)? din10 : din11;
assign mux_1_6 = (sel[0] == 0)? din12 : din13;
assign mux_1_7 = (sel[0] == 0)? din14 : din15;
assign mux_1_8 = (sel[0] == 0)? din16 : din17;
assign mux_1_9 = (sel[0] == 0)? din18 : din19;
assign mux_1_10 = (sel[0] == 0)? din20 : din21;
assign mux_1_11 = (sel[0] == 0)? din22 : din23;
assign mux_1_12 = (sel[0] == 0)? din24 : din25;
assign mux_1_13 = (sel[0] == 0)? din26 : din27;
assign mux_1_14 = (sel[0] == 0)? din28 : din29;
assign mux_1_15 = (sel[0] == 0)? din30 : din31;
assign mux_1_16 = (sel[0] == 0)? din32 : din33;
assign mux_1_17 = (sel[0] == 0)? din34 : din35;
assign mux_1_18 = (sel[0] == 0)? din36 : din37;
assign mux_1_19 = (sel[0] == 0)? din38 : din39;
assign mux_1_20 = (sel[0] == 0)? din40 : din41;
assign mux_1_21 = (sel[0] == 0)? din42 : din43;
assign mux_1_22 = (sel[0] == 0)? din44 : din45;
assign mux_1_23 = (sel[0] == 0)? din46 : din47;
assign mux_1_24 = (sel[0] == 0)? din48 : din49;
assign mux_1_25 = (sel[0] == 0)? din50 : din51;
assign mux_1_26 = (sel[0] == 0)? din52 : din53;
assign mux_1_27 = (sel[0] == 0)? din54 : din55;
assign mux_1_28 = (sel[0] == 0)? din56 : din57;
assign mux_1_29 = (sel[0] == 0)? din58 : din59;
assign mux_1_30 = (sel[0] == 0)? din60 : din61;
assign mux_1_31 = (sel[0] == 0)? din62 : din63;
assign mux_1_32 = (sel[0] == 0)? din64 : din65;
assign mux_1_33 = (sel[0] == 0)? din66 : din67;
assign mux_1_34 = (sel[0] == 0)? din68 : din69;
assign mux_1_35 = (sel[0] == 0)? din70 : din71;
assign mux_1_36 = (sel[0] == 0)? din72 : din73;
assign mux_1_37 = (sel[0] == 0)? din74 : din75;
assign mux_1_38 = (sel[0] == 0)? din76 : din77;
assign mux_1_39 = (sel[0] == 0)? din78 : din79;
assign mux_1_40 = (sel[0] == 0)? din80 : din81;
assign mux_1_41 = (sel[0] == 0)? din82 : din83;
assign mux_1_42 = (sel[0] == 0)? din84 : din85;
assign mux_1_43 = (sel[0] == 0)? din86 : din87;
assign mux_1_44 = (sel[0] == 0)? din88 : din89;
assign mux_1_45 = (sel[0] == 0)? din90 : din91;
assign mux_1_46 = (sel[0] == 0)? din92 : din93;
assign mux_1_47 = (sel[0] == 0)? din94 : din95;
assign mux_1_48 = (sel[0] == 0)? din96 : din97;
assign mux_1_49 = (sel[0] == 0)? din98 : din99;
assign mux_1_50 = (sel[0] == 0)? din100 : din101;
assign mux_1_51 = (sel[0] == 0)? din102 : din103;
assign mux_1_52 = (sel[0] == 0)? din104 : din105;
assign mux_1_53 = (sel[0] == 0)? din106 : din107;
assign mux_1_54 = (sel[0] == 0)? din108 : din109;
assign mux_1_55 = (sel[0] == 0)? din110 : din111;
assign mux_1_56 = (sel[0] == 0)? din112 : din113;
assign mux_1_57 = (sel[0] == 0)? din114 : din115;
assign mux_1_58 = (sel[0] == 0)? din116 : din117;
assign mux_1_59 = (sel[0] == 0)? din118 : din119;
assign mux_1_60 = (sel[0] == 0)? din120 : din121;
assign mux_1_61 = (sel[0] == 0)? din122 : din123;
assign mux_1_62 = (sel[0] == 0)? din124 : din125;
assign mux_1_63 = (sel[0] == 0)? din126 : din127;
assign mux_1_64 = (sel[0] == 0)? din128 : din129;
assign mux_1_65 = (sel[0] == 0)? din130 : din131;
assign mux_1_66 = (sel[0] == 0)? din132 : din133;
assign mux_1_67 = (sel[0] == 0)? din134 : din135;
assign mux_1_68 = (sel[0] == 0)? din136 : din137;
assign mux_1_69 = (sel[0] == 0)? din138 : din139;
assign mux_1_70 = (sel[0] == 0)? din140 : din141;
assign mux_1_71 = (sel[0] == 0)? din142 : din143;
assign mux_1_72 = (sel[0] == 0)? din144 : din145;
assign mux_1_73 = (sel[0] == 0)? din146 : din147;
assign mux_1_74 = (sel[0] == 0)? din148 : din149;
assign mux_1_75 = (sel[0] == 0)? din150 : din151;
assign mux_1_76 = (sel[0] == 0)? din152 : din153;
assign mux_1_77 = (sel[0] == 0)? din154 : din155;
assign mux_1_78 = (sel[0] == 0)? din156 : din157;
assign mux_1_79 = (sel[0] == 0)? din158 : din159;
assign mux_1_80 = (sel[0] == 0)? din160 : din161;
assign mux_1_81 = (sel[0] == 0)? din162 : din163;
assign mux_1_82 = (sel[0] == 0)? din164 : din165;
assign mux_1_83 = (sel[0] == 0)? din166 : din167;
assign mux_1_84 = (sel[0] == 0)? din168 : din169;
assign mux_1_85 = (sel[0] == 0)? din170 : din171;
assign mux_1_86 = (sel[0] == 0)? din172 : din173;
assign mux_1_87 = (sel[0] == 0)? din174 : din175;
assign mux_1_88 = (sel[0] == 0)? din176 : din177;
assign mux_1_89 = (sel[0] == 0)? din178 : din179;
assign mux_1_90 = (sel[0] == 0)? din180 : din181;
assign mux_1_91 = (sel[0] == 0)? din182 : din183;
assign mux_1_92 = (sel[0] == 0)? din184 : din185;
assign mux_1_93 = (sel[0] == 0)? din186 : din187;
assign mux_1_94 = (sel[0] == 0)? din188 : din189;
assign mux_1_95 = (sel[0] == 0)? din190 : din191;
assign mux_1_96 = (sel[0] == 0)? din192 : din193;
assign mux_1_97 = (sel[0] == 0)? din194 : din195;
assign mux_1_98 = (sel[0] == 0)? din196 : din197;
assign mux_1_99 = (sel[0] == 0)? din198 : din199;
assign mux_1_100 = (sel[0] == 0)? din200 : din201;
assign mux_1_101 = (sel[0] == 0)? din202 : din203;
assign mux_1_102 = (sel[0] == 0)? din204 : din205;
assign mux_1_103 = (sel[0] == 0)? din206 : din207;
assign mux_1_104 = (sel[0] == 0)? din208 : din209;
assign mux_1_105 = (sel[0] == 0)? din210 : din211;
assign mux_1_106 = (sel[0] == 0)? din212 : din213;
assign mux_1_107 = (sel[0] == 0)? din214 : din215;
assign mux_1_108 = (sel[0] == 0)? din216 : din217;
assign mux_1_109 = (sel[0] == 0)? din218 : din219;
assign mux_1_110 = (sel[0] == 0)? din220 : din221;
assign mux_1_111 = (sel[0] == 0)? din222 : din223;
assign mux_1_112 = (sel[0] == 0)? din224 : din225;
assign mux_1_113 = (sel[0] == 0)? din226 : din227;
assign mux_1_114 = (sel[0] == 0)? din228 : din229;
assign mux_1_115 = (sel[0] == 0)? din230 : din231;
assign mux_1_116 = (sel[0] == 0)? din232 : din233;
assign mux_1_117 = (sel[0] == 0)? din234 : din235;
assign mux_1_118 = (sel[0] == 0)? din236 : din237;
assign mux_1_119 = (sel[0] == 0)? din238 : din239;
assign mux_1_120 = (sel[0] == 0)? din240 : din241;
assign mux_1_121 = (sel[0] == 0)? din242 : din243;
assign mux_1_122 = (sel[0] == 0)? din244 : din245;
assign mux_1_123 = (sel[0] == 0)? din246 : din247;
assign mux_1_124 = (sel[0] == 0)? din248 : din249;
assign mux_1_125 = (sel[0] == 0)? din250 : din251;
assign mux_1_126 = (sel[0] == 0)? din252 : din253;
assign mux_1_127 = (sel[0] == 0)? din254 : din255;
assign mux_1_128 = (sel[0] == 0)? din256 : din257;
assign mux_1_129 = (sel[0] == 0)? din258 : din259;
assign mux_1_130 = (sel[0] == 0)? din260 : din261;
assign mux_1_131 = (sel[0] == 0)? din262 : din263;
assign mux_1_132 = (sel[0] == 0)? din264 : din265;
assign mux_1_133 = (sel[0] == 0)? din266 : din267;
assign mux_1_134 = (sel[0] == 0)? din268 : din269;
assign mux_1_135 = (sel[0] == 0)? din270 : din271;
assign mux_1_136 = (sel[0] == 0)? din272 : din273;
assign mux_1_137 = (sel[0] == 0)? din274 : din275;
assign mux_1_138 = (sel[0] == 0)? din276 : din277;
assign mux_1_139 = (sel[0] == 0)? din278 : din279;
assign mux_1_140 = (sel[0] == 0)? din280 : din281;
assign mux_1_141 = (sel[0] == 0)? din282 : din283;
assign mux_1_142 = (sel[0] == 0)? din284 : din285;
assign mux_1_143 = (sel[0] == 0)? din286 : din287;
assign mux_1_144 = (sel[0] == 0)? din288 : din289;
assign mux_1_145 = (sel[0] == 0)? din290 : din291;
assign mux_1_146 = (sel[0] == 0)? din292 : din293;
assign mux_1_147 = (sel[0] == 0)? din294 : din295;
assign mux_1_148 = (sel[0] == 0)? din296 : din297;
assign mux_1_149 = (sel[0] == 0)? din298 : din299;
assign mux_1_150 = (sel[0] == 0)? din300 : din301;
assign mux_1_151 = (sel[0] == 0)? din302 : din303;
assign mux_1_152 = (sel[0] == 0)? din304 : din305;
assign mux_1_153 = (sel[0] == 0)? din306 : din307;
assign mux_1_154 = (sel[0] == 0)? din308 : din309;
assign mux_1_155 = (sel[0] == 0)? din310 : din311;
assign mux_1_156 = (sel[0] == 0)? din312 : din313;
assign mux_1_157 = (sel[0] == 0)? din314 : din315;
assign mux_1_158 = (sel[0] == 0)? din316 : din317;
assign mux_1_159 = (sel[0] == 0)? din318 : din319;
assign mux_1_160 = (sel[0] == 0)? din320 : din321;
assign mux_1_161 = (sel[0] == 0)? din322 : din323;
assign mux_1_162 = (sel[0] == 0)? din324 : din325;
assign mux_1_163 = (sel[0] == 0)? din326 : din327;
assign mux_1_164 = (sel[0] == 0)? din328 : din329;
assign mux_1_165 = (sel[0] == 0)? din330 : din331;
assign mux_1_166 = (sel[0] == 0)? din332 : din333;
assign mux_1_167 = (sel[0] == 0)? din334 : din335;
assign mux_1_168 = (sel[0] == 0)? din336 : din337;
assign mux_1_169 = (sel[0] == 0)? din338 : din339;
assign mux_1_170 = (sel[0] == 0)? din340 : din341;
assign mux_1_171 = (sel[0] == 0)? din342 : din343;
assign mux_1_172 = (sel[0] == 0)? din344 : din345;
assign mux_1_173 = (sel[0] == 0)? din346 : din347;
assign mux_1_174 = (sel[0] == 0)? din348 : din349;
assign mux_1_175 = (sel[0] == 0)? din350 : din351;
assign mux_1_176 = (sel[0] == 0)? din352 : din353;
assign mux_1_177 = (sel[0] == 0)? din354 : din355;
assign mux_1_178 = (sel[0] == 0)? din356 : din357;
assign mux_1_179 = (sel[0] == 0)? din358 : din359;
assign mux_1_180 = (sel[0] == 0)? din360 : din361;
assign mux_1_181 = (sel[0] == 0)? din362 : din363;
assign mux_1_182 = (sel[0] == 0)? din364 : din365;
assign mux_1_183 = (sel[0] == 0)? din366 : din367;
assign mux_1_184 = (sel[0] == 0)? din368 : din369;
assign mux_1_185 = (sel[0] == 0)? din370 : din371;
assign mux_1_186 = (sel[0] == 0)? din372 : din373;
assign mux_1_187 = (sel[0] == 0)? din374 : din375;
assign mux_1_188 = (sel[0] == 0)? din376 : din377;
assign mux_1_189 = (sel[0] == 0)? din378 : din379;
assign mux_1_190 = (sel[0] == 0)? din380 : din381;
assign mux_1_191 = (sel[0] == 0)? din382 : din383;
assign mux_1_192 = (sel[0] == 0)? din384 : din385;
assign mux_1_193 = (sel[0] == 0)? din386 : din387;
assign mux_1_194 = (sel[0] == 0)? din388 : din389;
assign mux_1_195 = (sel[0] == 0)? din390 : din391;
assign mux_1_196 = (sel[0] == 0)? din392 : din393;
assign mux_1_197 = (sel[0] == 0)? din394 : din395;
assign mux_1_198 = (sel[0] == 0)? din396 : din397;
assign mux_1_199 = (sel[0] == 0)? din398 : din399;
assign mux_1_200 = (sel[0] == 0)? din400 : din401;
assign mux_1_201 = (sel[0] == 0)? din402 : din403;
assign mux_1_202 = (sel[0] == 0)? din404 : din405;
assign mux_1_203 = (sel[0] == 0)? din406 : din407;
assign mux_1_204 = (sel[0] == 0)? din408 : din409;
assign mux_1_205 = (sel[0] == 0)? din410 : din411;
assign mux_1_206 = (sel[0] == 0)? din412 : din413;
assign mux_1_207 = (sel[0] == 0)? din414 : din415;
assign mux_1_208 = (sel[0] == 0)? din416 : din417;
assign mux_1_209 = (sel[0] == 0)? din418 : din419;
assign mux_1_210 = (sel[0] == 0)? din420 : din421;
assign mux_1_211 = (sel[0] == 0)? din422 : din423;
assign mux_1_212 = (sel[0] == 0)? din424 : din425;
assign mux_1_213 = (sel[0] == 0)? din426 : din427;
assign mux_1_214 = (sel[0] == 0)? din428 : din429;
assign mux_1_215 = (sel[0] == 0)? din430 : din431;
assign mux_1_216 = (sel[0] == 0)? din432 : din433;
assign mux_1_217 = (sel[0] == 0)? din434 : din435;
assign mux_1_218 = (sel[0] == 0)? din436 : din437;
assign mux_1_219 = (sel[0] == 0)? din438 : din439;
assign mux_1_220 = (sel[0] == 0)? din440 : din441;
assign mux_1_221 = (sel[0] == 0)? din442 : din443;
assign mux_1_222 = (sel[0] == 0)? din444 : din445;
assign mux_1_223 = (sel[0] == 0)? din446 : din447;
assign mux_1_224 = (sel[0] == 0)? din448 : din449;
assign mux_1_225 = (sel[0] == 0)? din450 : din451;
assign mux_1_226 = (sel[0] == 0)? din452 : din453;
assign mux_1_227 = (sel[0] == 0)? din454 : din455;
assign mux_1_228 = (sel[0] == 0)? din456 : din457;
assign mux_1_229 = (sel[0] == 0)? din458 : din459;
assign mux_1_230 = (sel[0] == 0)? din460 : din461;
assign mux_1_231 = (sel[0] == 0)? din462 : din463;
assign mux_1_232 = (sel[0] == 0)? din464 : din465;
assign mux_1_233 = (sel[0] == 0)? din466 : din467;
assign mux_1_234 = (sel[0] == 0)? din468 : din469;
assign mux_1_235 = (sel[0] == 0)? din470 : din471;
assign mux_1_236 = (sel[0] == 0)? din472 : din473;
assign mux_1_237 = (sel[0] == 0)? din474 : din475;
assign mux_1_238 = (sel[0] == 0)? din476 : din477;
assign mux_1_239 = (sel[0] == 0)? din478 : din479;
assign mux_1_240 = (sel[0] == 0)? din480 : din481;
assign mux_1_241 = (sel[0] == 0)? din482 : din483;
assign mux_1_242 = (sel[0] == 0)? din484 : din485;
assign mux_1_243 = (sel[0] == 0)? din486 : din487;
assign mux_1_244 = (sel[0] == 0)? din488 : din489;
assign mux_1_245 = (sel[0] == 0)? din490 : din491;
assign mux_1_246 = (sel[0] == 0)? din492 : din493;
assign mux_1_247 = (sel[0] == 0)? din494 : din495;
assign mux_1_248 = (sel[0] == 0)? din496 : din497;
assign mux_1_249 = (sel[0] == 0)? din498 : din499;
assign mux_1_250 = (sel[0] == 0)? din500 : din501;
assign mux_1_251 = (sel[0] == 0)? din502 : din503;
assign mux_1_252 = (sel[0] == 0)? din504 : din505;
assign mux_1_253 = (sel[0] == 0)? din506 : din507;
assign mux_1_254 = (sel[0] == 0)? din508 : din509;
assign mux_1_255 = (sel[0] == 0)? din510 : din511;
assign mux_1_256 = (sel[0] == 0)? din512 : din513;
assign mux_1_257 = (sel[0] == 0)? din514 : din515;
assign mux_1_258 = (sel[0] == 0)? din516 : din517;
assign mux_1_259 = (sel[0] == 0)? din518 : din519;
assign mux_1_260 = (sel[0] == 0)? din520 : din521;
assign mux_1_261 = (sel[0] == 0)? din522 : din523;
assign mux_1_262 = (sel[0] == 0)? din524 : din525;
assign mux_1_263 = (sel[0] == 0)? din526 : din527;
assign mux_1_264 = (sel[0] == 0)? din528 : din529;
assign mux_1_265 = (sel[0] == 0)? din530 : din531;
assign mux_1_266 = (sel[0] == 0)? din532 : din533;
assign mux_1_267 = (sel[0] == 0)? din534 : din535;
assign mux_1_268 = (sel[0] == 0)? din536 : din537;
assign mux_1_269 = (sel[0] == 0)? din538 : din539;
assign mux_1_270 = (sel[0] == 0)? din540 : din541;
assign mux_1_271 = (sel[0] == 0)? din542 : din543;
assign mux_1_272 = (sel[0] == 0)? din544 : din545;
assign mux_1_273 = (sel[0] == 0)? din546 : din547;
assign mux_1_274 = (sel[0] == 0)? din548 : din549;
assign mux_1_275 = (sel[0] == 0)? din550 : din551;
assign mux_1_276 = (sel[0] == 0)? din552 : din553;
assign mux_1_277 = (sel[0] == 0)? din554 : din555;
assign mux_1_278 = (sel[0] == 0)? din556 : din557;
assign mux_1_279 = (sel[0] == 0)? din558 : din559;
assign mux_1_280 = (sel[0] == 0)? din560 : din561;
assign mux_1_281 = (sel[0] == 0)? din562 : din563;
assign mux_1_282 = (sel[0] == 0)? din564 : din565;
assign mux_1_283 = (sel[0] == 0)? din566 : din567;
assign mux_1_284 = (sel[0] == 0)? din568 : din569;
assign mux_1_285 = (sel[0] == 0)? din570 : din571;
assign mux_1_286 = (sel[0] == 0)? din572 : din573;
assign mux_1_287 = (sel[0] == 0)? din574 : din575;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;
assign mux_2_1 = (sel[1] == 0)? mux_1_2 : mux_1_3;
assign mux_2_2 = (sel[1] == 0)? mux_1_4 : mux_1_5;
assign mux_2_3 = (sel[1] == 0)? mux_1_6 : mux_1_7;
assign mux_2_4 = (sel[1] == 0)? mux_1_8 : mux_1_9;
assign mux_2_5 = (sel[1] == 0)? mux_1_10 : mux_1_11;
assign mux_2_6 = (sel[1] == 0)? mux_1_12 : mux_1_13;
assign mux_2_7 = (sel[1] == 0)? mux_1_14 : mux_1_15;
assign mux_2_8 = (sel[1] == 0)? mux_1_16 : mux_1_17;
assign mux_2_9 = (sel[1] == 0)? mux_1_18 : mux_1_19;
assign mux_2_10 = (sel[1] == 0)? mux_1_20 : mux_1_21;
assign mux_2_11 = (sel[1] == 0)? mux_1_22 : mux_1_23;
assign mux_2_12 = (sel[1] == 0)? mux_1_24 : mux_1_25;
assign mux_2_13 = (sel[1] == 0)? mux_1_26 : mux_1_27;
assign mux_2_14 = (sel[1] == 0)? mux_1_28 : mux_1_29;
assign mux_2_15 = (sel[1] == 0)? mux_1_30 : mux_1_31;
assign mux_2_16 = (sel[1] == 0)? mux_1_32 : mux_1_33;
assign mux_2_17 = (sel[1] == 0)? mux_1_34 : mux_1_35;
assign mux_2_18 = (sel[1] == 0)? mux_1_36 : mux_1_37;
assign mux_2_19 = (sel[1] == 0)? mux_1_38 : mux_1_39;
assign mux_2_20 = (sel[1] == 0)? mux_1_40 : mux_1_41;
assign mux_2_21 = (sel[1] == 0)? mux_1_42 : mux_1_43;
assign mux_2_22 = (sel[1] == 0)? mux_1_44 : mux_1_45;
assign mux_2_23 = (sel[1] == 0)? mux_1_46 : mux_1_47;
assign mux_2_24 = (sel[1] == 0)? mux_1_48 : mux_1_49;
assign mux_2_25 = (sel[1] == 0)? mux_1_50 : mux_1_51;
assign mux_2_26 = (sel[1] == 0)? mux_1_52 : mux_1_53;
assign mux_2_27 = (sel[1] == 0)? mux_1_54 : mux_1_55;
assign mux_2_28 = (sel[1] == 0)? mux_1_56 : mux_1_57;
assign mux_2_29 = (sel[1] == 0)? mux_1_58 : mux_1_59;
assign mux_2_30 = (sel[1] == 0)? mux_1_60 : mux_1_61;
assign mux_2_31 = (sel[1] == 0)? mux_1_62 : mux_1_63;
assign mux_2_32 = (sel[1] == 0)? mux_1_64 : mux_1_65;
assign mux_2_33 = (sel[1] == 0)? mux_1_66 : mux_1_67;
assign mux_2_34 = (sel[1] == 0)? mux_1_68 : mux_1_69;
assign mux_2_35 = (sel[1] == 0)? mux_1_70 : mux_1_71;
assign mux_2_36 = (sel[1] == 0)? mux_1_72 : mux_1_73;
assign mux_2_37 = (sel[1] == 0)? mux_1_74 : mux_1_75;
assign mux_2_38 = (sel[1] == 0)? mux_1_76 : mux_1_77;
assign mux_2_39 = (sel[1] == 0)? mux_1_78 : mux_1_79;
assign mux_2_40 = (sel[1] == 0)? mux_1_80 : mux_1_81;
assign mux_2_41 = (sel[1] == 0)? mux_1_82 : mux_1_83;
assign mux_2_42 = (sel[1] == 0)? mux_1_84 : mux_1_85;
assign mux_2_43 = (sel[1] == 0)? mux_1_86 : mux_1_87;
assign mux_2_44 = (sel[1] == 0)? mux_1_88 : mux_1_89;
assign mux_2_45 = (sel[1] == 0)? mux_1_90 : mux_1_91;
assign mux_2_46 = (sel[1] == 0)? mux_1_92 : mux_1_93;
assign mux_2_47 = (sel[1] == 0)? mux_1_94 : mux_1_95;
assign mux_2_48 = (sel[1] == 0)? mux_1_96 : mux_1_97;
assign mux_2_49 = (sel[1] == 0)? mux_1_98 : mux_1_99;
assign mux_2_50 = (sel[1] == 0)? mux_1_100 : mux_1_101;
assign mux_2_51 = (sel[1] == 0)? mux_1_102 : mux_1_103;
assign mux_2_52 = (sel[1] == 0)? mux_1_104 : mux_1_105;
assign mux_2_53 = (sel[1] == 0)? mux_1_106 : mux_1_107;
assign mux_2_54 = (sel[1] == 0)? mux_1_108 : mux_1_109;
assign mux_2_55 = (sel[1] == 0)? mux_1_110 : mux_1_111;
assign mux_2_56 = (sel[1] == 0)? mux_1_112 : mux_1_113;
assign mux_2_57 = (sel[1] == 0)? mux_1_114 : mux_1_115;
assign mux_2_58 = (sel[1] == 0)? mux_1_116 : mux_1_117;
assign mux_2_59 = (sel[1] == 0)? mux_1_118 : mux_1_119;
assign mux_2_60 = (sel[1] == 0)? mux_1_120 : mux_1_121;
assign mux_2_61 = (sel[1] == 0)? mux_1_122 : mux_1_123;
assign mux_2_62 = (sel[1] == 0)? mux_1_124 : mux_1_125;
assign mux_2_63 = (sel[1] == 0)? mux_1_126 : mux_1_127;
assign mux_2_64 = (sel[1] == 0)? mux_1_128 : mux_1_129;
assign mux_2_65 = (sel[1] == 0)? mux_1_130 : mux_1_131;
assign mux_2_66 = (sel[1] == 0)? mux_1_132 : mux_1_133;
assign mux_2_67 = (sel[1] == 0)? mux_1_134 : mux_1_135;
assign mux_2_68 = (sel[1] == 0)? mux_1_136 : mux_1_137;
assign mux_2_69 = (sel[1] == 0)? mux_1_138 : mux_1_139;
assign mux_2_70 = (sel[1] == 0)? mux_1_140 : mux_1_141;
assign mux_2_71 = (sel[1] == 0)? mux_1_142 : mux_1_143;
assign mux_2_72 = (sel[1] == 0)? mux_1_144 : mux_1_145;
assign mux_2_73 = (sel[1] == 0)? mux_1_146 : mux_1_147;
assign mux_2_74 = (sel[1] == 0)? mux_1_148 : mux_1_149;
assign mux_2_75 = (sel[1] == 0)? mux_1_150 : mux_1_151;
assign mux_2_76 = (sel[1] == 0)? mux_1_152 : mux_1_153;
assign mux_2_77 = (sel[1] == 0)? mux_1_154 : mux_1_155;
assign mux_2_78 = (sel[1] == 0)? mux_1_156 : mux_1_157;
assign mux_2_79 = (sel[1] == 0)? mux_1_158 : mux_1_159;
assign mux_2_80 = (sel[1] == 0)? mux_1_160 : mux_1_161;
assign mux_2_81 = (sel[1] == 0)? mux_1_162 : mux_1_163;
assign mux_2_82 = (sel[1] == 0)? mux_1_164 : mux_1_165;
assign mux_2_83 = (sel[1] == 0)? mux_1_166 : mux_1_167;
assign mux_2_84 = (sel[1] == 0)? mux_1_168 : mux_1_169;
assign mux_2_85 = (sel[1] == 0)? mux_1_170 : mux_1_171;
assign mux_2_86 = (sel[1] == 0)? mux_1_172 : mux_1_173;
assign mux_2_87 = (sel[1] == 0)? mux_1_174 : mux_1_175;
assign mux_2_88 = (sel[1] == 0)? mux_1_176 : mux_1_177;
assign mux_2_89 = (sel[1] == 0)? mux_1_178 : mux_1_179;
assign mux_2_90 = (sel[1] == 0)? mux_1_180 : mux_1_181;
assign mux_2_91 = (sel[1] == 0)? mux_1_182 : mux_1_183;
assign mux_2_92 = (sel[1] == 0)? mux_1_184 : mux_1_185;
assign mux_2_93 = (sel[1] == 0)? mux_1_186 : mux_1_187;
assign mux_2_94 = (sel[1] == 0)? mux_1_188 : mux_1_189;
assign mux_2_95 = (sel[1] == 0)? mux_1_190 : mux_1_191;
assign mux_2_96 = (sel[1] == 0)? mux_1_192 : mux_1_193;
assign mux_2_97 = (sel[1] == 0)? mux_1_194 : mux_1_195;
assign mux_2_98 = (sel[1] == 0)? mux_1_196 : mux_1_197;
assign mux_2_99 = (sel[1] == 0)? mux_1_198 : mux_1_199;
assign mux_2_100 = (sel[1] == 0)? mux_1_200 : mux_1_201;
assign mux_2_101 = (sel[1] == 0)? mux_1_202 : mux_1_203;
assign mux_2_102 = (sel[1] == 0)? mux_1_204 : mux_1_205;
assign mux_2_103 = (sel[1] == 0)? mux_1_206 : mux_1_207;
assign mux_2_104 = (sel[1] == 0)? mux_1_208 : mux_1_209;
assign mux_2_105 = (sel[1] == 0)? mux_1_210 : mux_1_211;
assign mux_2_106 = (sel[1] == 0)? mux_1_212 : mux_1_213;
assign mux_2_107 = (sel[1] == 0)? mux_1_214 : mux_1_215;
assign mux_2_108 = (sel[1] == 0)? mux_1_216 : mux_1_217;
assign mux_2_109 = (sel[1] == 0)? mux_1_218 : mux_1_219;
assign mux_2_110 = (sel[1] == 0)? mux_1_220 : mux_1_221;
assign mux_2_111 = (sel[1] == 0)? mux_1_222 : mux_1_223;
assign mux_2_112 = (sel[1] == 0)? mux_1_224 : mux_1_225;
assign mux_2_113 = (sel[1] == 0)? mux_1_226 : mux_1_227;
assign mux_2_114 = (sel[1] == 0)? mux_1_228 : mux_1_229;
assign mux_2_115 = (sel[1] == 0)? mux_1_230 : mux_1_231;
assign mux_2_116 = (sel[1] == 0)? mux_1_232 : mux_1_233;
assign mux_2_117 = (sel[1] == 0)? mux_1_234 : mux_1_235;
assign mux_2_118 = (sel[1] == 0)? mux_1_236 : mux_1_237;
assign mux_2_119 = (sel[1] == 0)? mux_1_238 : mux_1_239;
assign mux_2_120 = (sel[1] == 0)? mux_1_240 : mux_1_241;
assign mux_2_121 = (sel[1] == 0)? mux_1_242 : mux_1_243;
assign mux_2_122 = (sel[1] == 0)? mux_1_244 : mux_1_245;
assign mux_2_123 = (sel[1] == 0)? mux_1_246 : mux_1_247;
assign mux_2_124 = (sel[1] == 0)? mux_1_248 : mux_1_249;
assign mux_2_125 = (sel[1] == 0)? mux_1_250 : mux_1_251;
assign mux_2_126 = (sel[1] == 0)? mux_1_252 : mux_1_253;
assign mux_2_127 = (sel[1] == 0)? mux_1_254 : mux_1_255;
assign mux_2_128 = (sel[1] == 0)? mux_1_256 : mux_1_257;
assign mux_2_129 = (sel[1] == 0)? mux_1_258 : mux_1_259;
assign mux_2_130 = (sel[1] == 0)? mux_1_260 : mux_1_261;
assign mux_2_131 = (sel[1] == 0)? mux_1_262 : mux_1_263;
assign mux_2_132 = (sel[1] == 0)? mux_1_264 : mux_1_265;
assign mux_2_133 = (sel[1] == 0)? mux_1_266 : mux_1_267;
assign mux_2_134 = (sel[1] == 0)? mux_1_268 : mux_1_269;
assign mux_2_135 = (sel[1] == 0)? mux_1_270 : mux_1_271;
assign mux_2_136 = (sel[1] == 0)? mux_1_272 : mux_1_273;
assign mux_2_137 = (sel[1] == 0)? mux_1_274 : mux_1_275;
assign mux_2_138 = (sel[1] == 0)? mux_1_276 : mux_1_277;
assign mux_2_139 = (sel[1] == 0)? mux_1_278 : mux_1_279;
assign mux_2_140 = (sel[1] == 0)? mux_1_280 : mux_1_281;
assign mux_2_141 = (sel[1] == 0)? mux_1_282 : mux_1_283;
assign mux_2_142 = (sel[1] == 0)? mux_1_284 : mux_1_285;
assign mux_2_143 = (sel[1] == 0)? mux_1_286 : mux_1_287;

// Generate level 3 logic
assign mux_3_0 = (sel[2] == 0)? mux_2_0 : mux_2_1;
assign mux_3_1 = (sel[2] == 0)? mux_2_2 : mux_2_3;
assign mux_3_2 = (sel[2] == 0)? mux_2_4 : mux_2_5;
assign mux_3_3 = (sel[2] == 0)? mux_2_6 : mux_2_7;
assign mux_3_4 = (sel[2] == 0)? mux_2_8 : mux_2_9;
assign mux_3_5 = (sel[2] == 0)? mux_2_10 : mux_2_11;
assign mux_3_6 = (sel[2] == 0)? mux_2_12 : mux_2_13;
assign mux_3_7 = (sel[2] == 0)? mux_2_14 : mux_2_15;
assign mux_3_8 = (sel[2] == 0)? mux_2_16 : mux_2_17;
assign mux_3_9 = (sel[2] == 0)? mux_2_18 : mux_2_19;
assign mux_3_10 = (sel[2] == 0)? mux_2_20 : mux_2_21;
assign mux_3_11 = (sel[2] == 0)? mux_2_22 : mux_2_23;
assign mux_3_12 = (sel[2] == 0)? mux_2_24 : mux_2_25;
assign mux_3_13 = (sel[2] == 0)? mux_2_26 : mux_2_27;
assign mux_3_14 = (sel[2] == 0)? mux_2_28 : mux_2_29;
assign mux_3_15 = (sel[2] == 0)? mux_2_30 : mux_2_31;
assign mux_3_16 = (sel[2] == 0)? mux_2_32 : mux_2_33;
assign mux_3_17 = (sel[2] == 0)? mux_2_34 : mux_2_35;
assign mux_3_18 = (sel[2] == 0)? mux_2_36 : mux_2_37;
assign mux_3_19 = (sel[2] == 0)? mux_2_38 : mux_2_39;
assign mux_3_20 = (sel[2] == 0)? mux_2_40 : mux_2_41;
assign mux_3_21 = (sel[2] == 0)? mux_2_42 : mux_2_43;
assign mux_3_22 = (sel[2] == 0)? mux_2_44 : mux_2_45;
assign mux_3_23 = (sel[2] == 0)? mux_2_46 : mux_2_47;
assign mux_3_24 = (sel[2] == 0)? mux_2_48 : mux_2_49;
assign mux_3_25 = (sel[2] == 0)? mux_2_50 : mux_2_51;
assign mux_3_26 = (sel[2] == 0)? mux_2_52 : mux_2_53;
assign mux_3_27 = (sel[2] == 0)? mux_2_54 : mux_2_55;
assign mux_3_28 = (sel[2] == 0)? mux_2_56 : mux_2_57;
assign mux_3_29 = (sel[2] == 0)? mux_2_58 : mux_2_59;
assign mux_3_30 = (sel[2] == 0)? mux_2_60 : mux_2_61;
assign mux_3_31 = (sel[2] == 0)? mux_2_62 : mux_2_63;
assign mux_3_32 = (sel[2] == 0)? mux_2_64 : mux_2_65;
assign mux_3_33 = (sel[2] == 0)? mux_2_66 : mux_2_67;
assign mux_3_34 = (sel[2] == 0)? mux_2_68 : mux_2_69;
assign mux_3_35 = (sel[2] == 0)? mux_2_70 : mux_2_71;
assign mux_3_36 = (sel[2] == 0)? mux_2_72 : mux_2_73;
assign mux_3_37 = (sel[2] == 0)? mux_2_74 : mux_2_75;
assign mux_3_38 = (sel[2] == 0)? mux_2_76 : mux_2_77;
assign mux_3_39 = (sel[2] == 0)? mux_2_78 : mux_2_79;
assign mux_3_40 = (sel[2] == 0)? mux_2_80 : mux_2_81;
assign mux_3_41 = (sel[2] == 0)? mux_2_82 : mux_2_83;
assign mux_3_42 = (sel[2] == 0)? mux_2_84 : mux_2_85;
assign mux_3_43 = (sel[2] == 0)? mux_2_86 : mux_2_87;
assign mux_3_44 = (sel[2] == 0)? mux_2_88 : mux_2_89;
assign mux_3_45 = (sel[2] == 0)? mux_2_90 : mux_2_91;
assign mux_3_46 = (sel[2] == 0)? mux_2_92 : mux_2_93;
assign mux_3_47 = (sel[2] == 0)? mux_2_94 : mux_2_95;
assign mux_3_48 = (sel[2] == 0)? mux_2_96 : mux_2_97;
assign mux_3_49 = (sel[2] == 0)? mux_2_98 : mux_2_99;
assign mux_3_50 = (sel[2] == 0)? mux_2_100 : mux_2_101;
assign mux_3_51 = (sel[2] == 0)? mux_2_102 : mux_2_103;
assign mux_3_52 = (sel[2] == 0)? mux_2_104 : mux_2_105;
assign mux_3_53 = (sel[2] == 0)? mux_2_106 : mux_2_107;
assign mux_3_54 = (sel[2] == 0)? mux_2_108 : mux_2_109;
assign mux_3_55 = (sel[2] == 0)? mux_2_110 : mux_2_111;
assign mux_3_56 = (sel[2] == 0)? mux_2_112 : mux_2_113;
assign mux_3_57 = (sel[2] == 0)? mux_2_114 : mux_2_115;
assign mux_3_58 = (sel[2] == 0)? mux_2_116 : mux_2_117;
assign mux_3_59 = (sel[2] == 0)? mux_2_118 : mux_2_119;
assign mux_3_60 = (sel[2] == 0)? mux_2_120 : mux_2_121;
assign mux_3_61 = (sel[2] == 0)? mux_2_122 : mux_2_123;
assign mux_3_62 = (sel[2] == 0)? mux_2_124 : mux_2_125;
assign mux_3_63 = (sel[2] == 0)? mux_2_126 : mux_2_127;
assign mux_3_64 = (sel[2] == 0)? mux_2_128 : mux_2_129;
assign mux_3_65 = (sel[2] == 0)? mux_2_130 : mux_2_131;
assign mux_3_66 = (sel[2] == 0)? mux_2_132 : mux_2_133;
assign mux_3_67 = (sel[2] == 0)? mux_2_134 : mux_2_135;
assign mux_3_68 = (sel[2] == 0)? mux_2_136 : mux_2_137;
assign mux_3_69 = (sel[2] == 0)? mux_2_138 : mux_2_139;
assign mux_3_70 = (sel[2] == 0)? mux_2_140 : mux_2_141;
assign mux_3_71 = (sel[2] == 0)? mux_2_142 : mux_2_143;

// Generate level 4 logic
assign mux_4_0 = (sel[3] == 0)? mux_3_0 : mux_3_1;
assign mux_4_1 = (sel[3] == 0)? mux_3_2 : mux_3_3;
assign mux_4_2 = (sel[3] == 0)? mux_3_4 : mux_3_5;
assign mux_4_3 = (sel[3] == 0)? mux_3_6 : mux_3_7;
assign mux_4_4 = (sel[3] == 0)? mux_3_8 : mux_3_9;
assign mux_4_5 = (sel[3] == 0)? mux_3_10 : mux_3_11;
assign mux_4_6 = (sel[3] == 0)? mux_3_12 : mux_3_13;
assign mux_4_7 = (sel[3] == 0)? mux_3_14 : mux_3_15;
assign mux_4_8 = (sel[3] == 0)? mux_3_16 : mux_3_17;
assign mux_4_9 = (sel[3] == 0)? mux_3_18 : mux_3_19;
assign mux_4_10 = (sel[3] == 0)? mux_3_20 : mux_3_21;
assign mux_4_11 = (sel[3] == 0)? mux_3_22 : mux_3_23;
assign mux_4_12 = (sel[3] == 0)? mux_3_24 : mux_3_25;
assign mux_4_13 = (sel[3] == 0)? mux_3_26 : mux_3_27;
assign mux_4_14 = (sel[3] == 0)? mux_3_28 : mux_3_29;
assign mux_4_15 = (sel[3] == 0)? mux_3_30 : mux_3_31;
assign mux_4_16 = (sel[3] == 0)? mux_3_32 : mux_3_33;
assign mux_4_17 = (sel[3] == 0)? mux_3_34 : mux_3_35;
assign mux_4_18 = (sel[3] == 0)? mux_3_36 : mux_3_37;
assign mux_4_19 = (sel[3] == 0)? mux_3_38 : mux_3_39;
assign mux_4_20 = (sel[3] == 0)? mux_3_40 : mux_3_41;
assign mux_4_21 = (sel[3] == 0)? mux_3_42 : mux_3_43;
assign mux_4_22 = (sel[3] == 0)? mux_3_44 : mux_3_45;
assign mux_4_23 = (sel[3] == 0)? mux_3_46 : mux_3_47;
assign mux_4_24 = (sel[3] == 0)? mux_3_48 : mux_3_49;
assign mux_4_25 = (sel[3] == 0)? mux_3_50 : mux_3_51;
assign mux_4_26 = (sel[3] == 0)? mux_3_52 : mux_3_53;
assign mux_4_27 = (sel[3] == 0)? mux_3_54 : mux_3_55;
assign mux_4_28 = (sel[3] == 0)? mux_3_56 : mux_3_57;
assign mux_4_29 = (sel[3] == 0)? mux_3_58 : mux_3_59;
assign mux_4_30 = (sel[3] == 0)? mux_3_60 : mux_3_61;
assign mux_4_31 = (sel[3] == 0)? mux_3_62 : mux_3_63;
assign mux_4_32 = (sel[3] == 0)? mux_3_64 : mux_3_65;
assign mux_4_33 = (sel[3] == 0)? mux_3_66 : mux_3_67;
assign mux_4_34 = (sel[3] == 0)? mux_3_68 : mux_3_69;
assign mux_4_35 = (sel[3] == 0)? mux_3_70 : mux_3_71;

// Generate level 5 logic
assign mux_5_0 = (sel[4] == 0)? mux_4_0 : mux_4_1;
assign mux_5_1 = (sel[4] == 0)? mux_4_2 : mux_4_3;
assign mux_5_2 = (sel[4] == 0)? mux_4_4 : mux_4_5;
assign mux_5_3 = (sel[4] == 0)? mux_4_6 : mux_4_7;
assign mux_5_4 = (sel[4] == 0)? mux_4_8 : mux_4_9;
assign mux_5_5 = (sel[4] == 0)? mux_4_10 : mux_4_11;
assign mux_5_6 = (sel[4] == 0)? mux_4_12 : mux_4_13;
assign mux_5_7 = (sel[4] == 0)? mux_4_14 : mux_4_15;
assign mux_5_8 = (sel[4] == 0)? mux_4_16 : mux_4_17;
assign mux_5_9 = (sel[4] == 0)? mux_4_18 : mux_4_19;
assign mux_5_10 = (sel[4] == 0)? mux_4_20 : mux_4_21;
assign mux_5_11 = (sel[4] == 0)? mux_4_22 : mux_4_23;
assign mux_5_12 = (sel[4] == 0)? mux_4_24 : mux_4_25;
assign mux_5_13 = (sel[4] == 0)? mux_4_26 : mux_4_27;
assign mux_5_14 = (sel[4] == 0)? mux_4_28 : mux_4_29;
assign mux_5_15 = (sel[4] == 0)? mux_4_30 : mux_4_31;
assign mux_5_16 = (sel[4] == 0)? mux_4_32 : mux_4_33;
assign mux_5_17 = (sel[4] == 0)? mux_4_34 : mux_4_35;

// Generate level 6 logic
assign mux_6_0 = (sel[5] == 0)? mux_5_0 : mux_5_1;
assign mux_6_1 = (sel[5] == 0)? mux_5_2 : mux_5_3;
assign mux_6_2 = (sel[5] == 0)? mux_5_4 : mux_5_5;
assign mux_6_3 = (sel[5] == 0)? mux_5_6 : mux_5_7;
assign mux_6_4 = (sel[5] == 0)? mux_5_8 : mux_5_9;
assign mux_6_5 = (sel[5] == 0)? mux_5_10 : mux_5_11;
assign mux_6_6 = (sel[5] == 0)? mux_5_12 : mux_5_13;
assign mux_6_7 = (sel[5] == 0)? mux_5_14 : mux_5_15;
assign mux_6_8 = (sel[5] == 0)? mux_5_16 : mux_5_17;

// Generate level 7 logic
assign mux_7_0 = (sel[6] == 0)? mux_6_0 : mux_6_1;
assign mux_7_1 = (sel[6] == 0)? mux_6_2 : mux_6_3;
assign mux_7_2 = (sel[6] == 0)? mux_6_4 : mux_6_5;
assign mux_7_3 = (sel[6] == 0)? mux_6_6 : mux_6_7;
assign mux_7_4 = mux_6_8;

// Generate level 8 logic
assign mux_8_0 = (sel[7] == 0)? mux_7_0 : mux_7_1;
assign mux_8_1 = (sel[7] == 0)? mux_7_2 : mux_7_3;
assign mux_8_2 = mux_7_4;

// Generate level 9 logic
assign mux_9_0 = (sel[8] == 0)? mux_8_0 : mux_8_1;
assign mux_9_1 = mux_8_2;

// Generate level 10 logic
assign mux_10_0 = (sel[9] == 0)? mux_9_0 : mux_9_1;

// output logic
assign dout = mux_10_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Act4jc.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Act4jc_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Act4jc_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Act4jc(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Act4jc_rom StreamingFCLayer_Batch_3_Matrix_Vector_Act4jc_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc8D.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcc8D_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc8D_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcc8D(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcc8D_rom Thresholding_Batch_0_Thresholding_Batcc8D_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Acthbi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Acthbi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Acthbi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Acthbi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Acthbi_rom StreamingFCLayer_Batch_3_Matrix_Vector_Acthbi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActkbM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActkbM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActkbM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActkbM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActkbM_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActkbM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcLf8.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcLf8_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcLf8_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcLf8(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcLf8_rom Thresholding_Batch_0_Thresholding_BatcLf8_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbwn.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbwn_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbwn_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbwn(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbwn_rom Thresholding_Batch_0_Thresholding_Batcbwn_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_14_0/synth/finn_design_StreamingFIFO_14_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_14:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_14,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_14_0,StreamingFIFO_14,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_14_0,StreamingFIFO_14,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_14,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_14_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_14 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_Batccud.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_Batccud_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_Batccud_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_Batccud(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_Batccud_rom Thresholding_Batch_1_Thresholding_Batccud_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_ConvolutionInputGenerator_2_0/synth/finn_design_ConvolutionInputGenerator_2_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:ConvolutionInputGenerator_2:1.0
// IP Revision: 2101301317

(* X_CORE_INFO = "ConvolutionInputGenerator_2_ConvolutionInputGenerator_2,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_ConvolutionInputGenerator_2_0,ConvolutionInputGenerator_2_ConvolutionInputGenerator_2,{}" *)
(* CORE_GENERATION_INFO = "finn_design_ConvolutionInputGenerator_2_0,ConvolutionInputGenerator_2_ConvolutionInputGenerator_2,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=ConvolutionInputGenerator_2,x_ipVersion=1.0,x_ipCoreRevision=2101301317,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_ConvolutionInputGenerator_2_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 3, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [23 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 3, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [23 : 0] out_V_V_TDATA;

  ConvolutionInputGenerator_2_ConvolutionInputGenerator_2 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Act3i2.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Act3i2_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Act3i2_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Act3i2(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Act3i2_rom StreamingFCLayer_Batch_2_Matrix_Vector_Act3i2_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batctde.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batctde_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 5;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batctde_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batctde(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd5;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batctde_rom Thresholding_Batch_0_Thresholding_Batctde_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcchv.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcchv_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcchv_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcchv(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcchv_rom Thresholding_Batch_0_Thresholding_Batcchv_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_0_0/synth/finn_design_StreamingFIFO_0_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_0:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_0,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_0_0,StreamingFIFO_0,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_0_0,StreamingFIFO_0,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_0,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_0_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [7 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_0 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Activa.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingFCLayer_Batch_2_Matrix_Vector_Activa (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY,
        weight_V_V_TDATA,
        weight_V_V_TVALID,
        weight_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state6 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [23:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;
input  [47:0] weight_V_V_TDATA;
input   weight_V_V_TVALID;
output   weight_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;
reg weight_V_V_TREADY;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] threshs_m_thresholds_55_address0;
reg    threshs_m_thresholds_55_ce0;
wire   [15:0] threshs_m_thresholds_55_q0;
wire   [3:0] threshs_m_thresholds_54_address0;
reg    threshs_m_thresholds_54_ce0;
wire   [15:0] threshs_m_thresholds_54_q0;
wire   [3:0] threshs_m_thresholds_49_address0;
reg    threshs_m_thresholds_49_ce0;
wire   [15:0] threshs_m_thresholds_49_q0;
wire   [3:0] threshs_m_thresholds_48_address0;
reg    threshs_m_thresholds_48_ce0;
wire   [15:0] threshs_m_thresholds_48_q0;
wire   [3:0] threshs_m_thresholds_47_address0;
reg    threshs_m_thresholds_47_ce0;
wire   [15:0] threshs_m_thresholds_47_q0;
wire   [3:0] threshs_m_thresholds_46_address0;
reg    threshs_m_thresholds_46_ce0;
wire   [15:0] threshs_m_thresholds_46_q0;
wire   [3:0] threshs_m_thresholds_45_address0;
reg    threshs_m_thresholds_45_ce0;
wire   [15:0] threshs_m_thresholds_45_q0;
wire   [3:0] threshs_m_thresholds_44_address0;
reg    threshs_m_thresholds_44_ce0;
wire   [15:0] threshs_m_thresholds_44_q0;
wire   [3:0] threshs_m_thresholds_43_address0;
reg    threshs_m_thresholds_43_ce0;
wire   [15:0] threshs_m_thresholds_43_q0;
wire   [3:0] threshs_m_thresholds_42_address0;
reg    threshs_m_thresholds_42_ce0;
wire   [15:0] threshs_m_thresholds_42_q0;
wire   [3:0] threshs_m_thresholds_53_address0;
reg    threshs_m_thresholds_53_ce0;
wire   [15:0] threshs_m_thresholds_53_q0;
wire   [3:0] threshs_m_thresholds_52_address0;
reg    threshs_m_thresholds_52_ce0;
wire   [15:0] threshs_m_thresholds_52_q0;
wire   [3:0] threshs_m_thresholds_51_address0;
reg    threshs_m_thresholds_51_ce0;
wire   [15:0] threshs_m_thresholds_51_q0;
wire   [3:0] threshs_m_thresholds_50_address0;
reg    threshs_m_thresholds_50_ce0;
wire   [15:0] threshs_m_thresholds_50_q0;
wire   [3:0] threshs_m_thresholds_41_address0;
reg    threshs_m_thresholds_41_ce0;
wire   [15:0] threshs_m_thresholds_41_q0;
wire   [3:0] threshs_m_thresholds_40_address0;
reg    threshs_m_thresholds_40_ce0;
wire   [15:0] threshs_m_thresholds_40_q0;
wire   [3:0] threshs_m_thresholds_35_address0;
reg    threshs_m_thresholds_35_ce0;
wire   [15:0] threshs_m_thresholds_35_q0;
wire   [3:0] threshs_m_thresholds_34_address0;
reg    threshs_m_thresholds_34_ce0;
wire   [15:0] threshs_m_thresholds_34_q0;
wire   [3:0] threshs_m_thresholds_33_address0;
reg    threshs_m_thresholds_33_ce0;
wire   [15:0] threshs_m_thresholds_33_q0;
wire   [3:0] threshs_m_thresholds_32_address0;
reg    threshs_m_thresholds_32_ce0;
wire   [15:0] threshs_m_thresholds_32_q0;
wire   [3:0] threshs_m_thresholds_31_address0;
reg    threshs_m_thresholds_31_ce0;
wire   [15:0] threshs_m_thresholds_31_q0;
wire   [3:0] threshs_m_thresholds_30_address0;
reg    threshs_m_thresholds_30_ce0;
wire   [15:0] threshs_m_thresholds_30_q0;
wire   [3:0] threshs_m_thresholds_29_address0;
reg    threshs_m_thresholds_29_ce0;
wire   [15:0] threshs_m_thresholds_29_q0;
wire   [3:0] threshs_m_thresholds_28_address0;
reg    threshs_m_thresholds_28_ce0;
wire   [15:0] threshs_m_thresholds_28_q0;
wire   [3:0] threshs_m_thresholds_39_address0;
reg    threshs_m_thresholds_39_ce0;
wire   [15:0] threshs_m_thresholds_39_q0;
wire   [3:0] threshs_m_thresholds_38_address0;
reg    threshs_m_thresholds_38_ce0;
wire   [15:0] threshs_m_thresholds_38_q0;
wire   [3:0] threshs_m_thresholds_37_address0;
reg    threshs_m_thresholds_37_ce0;
wire   [15:0] threshs_m_thresholds_37_q0;
wire   [3:0] threshs_m_thresholds_36_address0;
reg    threshs_m_thresholds_36_ce0;
wire   [15:0] threshs_m_thresholds_36_q0;
wire   [3:0] threshs_m_thresholds_27_address0;
reg    threshs_m_thresholds_27_ce0;
wire   [15:0] threshs_m_thresholds_27_q0;
wire   [3:0] threshs_m_thresholds_26_address0;
reg    threshs_m_thresholds_26_ce0;
wire   [15:0] threshs_m_thresholds_26_q0;
wire   [3:0] threshs_m_thresholds_21_address0;
reg    threshs_m_thresholds_21_ce0;
wire   [15:0] threshs_m_thresholds_21_q0;
wire   [3:0] threshs_m_thresholds_20_address0;
reg    threshs_m_thresholds_20_ce0;
wire   [15:0] threshs_m_thresholds_20_q0;
wire   [3:0] threshs_m_thresholds_19_address0;
reg    threshs_m_thresholds_19_ce0;
wire   [15:0] threshs_m_thresholds_19_q0;
wire   [3:0] threshs_m_thresholds_18_address0;
reg    threshs_m_thresholds_18_ce0;
wire   [15:0] threshs_m_thresholds_18_q0;
wire   [3:0] threshs_m_thresholds_17_address0;
reg    threshs_m_thresholds_17_ce0;
wire   [15:0] threshs_m_thresholds_17_q0;
wire   [3:0] threshs_m_thresholds_16_address0;
reg    threshs_m_thresholds_16_ce0;
wire   [15:0] threshs_m_thresholds_16_q0;
wire   [3:0] threshs_m_thresholds_15_address0;
reg    threshs_m_thresholds_15_ce0;
wire   [15:0] threshs_m_thresholds_15_q0;
wire   [3:0] threshs_m_thresholds_14_address0;
reg    threshs_m_thresholds_14_ce0;
wire   [15:0] threshs_m_thresholds_14_q0;
wire   [3:0] threshs_m_thresholds_25_address0;
reg    threshs_m_thresholds_25_ce0;
wire   [15:0] threshs_m_thresholds_25_q0;
wire   [3:0] threshs_m_thresholds_24_address0;
reg    threshs_m_thresholds_24_ce0;
wire   [15:0] threshs_m_thresholds_24_q0;
wire   [3:0] threshs_m_thresholds_23_address0;
reg    threshs_m_thresholds_23_ce0;
wire   [15:0] threshs_m_thresholds_23_q0;
wire   [3:0] threshs_m_thresholds_22_address0;
reg    threshs_m_thresholds_22_ce0;
wire   [15:0] threshs_m_thresholds_22_q0;
wire   [3:0] threshs_m_thresholds_13_address0;
reg    threshs_m_thresholds_13_ce0;
wire   [15:0] threshs_m_thresholds_13_q0;
wire   [3:0] threshs_m_thresholds_12_address0;
reg    threshs_m_thresholds_12_ce0;
wire   [15:0] threshs_m_thresholds_12_q0;
wire   [3:0] threshs_m_thresholds_7_address0;
reg    threshs_m_thresholds_7_ce0;
wire   [15:0] threshs_m_thresholds_7_q0;
wire   [3:0] threshs_m_thresholds_6_address0;
reg    threshs_m_thresholds_6_ce0;
wire   [15:0] threshs_m_thresholds_6_q0;
wire   [3:0] threshs_m_thresholds_5_address0;
reg    threshs_m_thresholds_5_ce0;
wire   [15:0] threshs_m_thresholds_5_q0;
wire   [3:0] threshs_m_thresholds_4_address0;
reg    threshs_m_thresholds_4_ce0;
wire   [15:0] threshs_m_thresholds_4_q0;
wire   [3:0] threshs_m_thresholds_3_address0;
reg    threshs_m_thresholds_3_ce0;
wire   [15:0] threshs_m_thresholds_3_q0;
wire   [3:0] threshs_m_thresholds_2_address0;
reg    threshs_m_thresholds_2_ce0;
wire   [15:0] threshs_m_thresholds_2_q0;
wire   [3:0] threshs_m_thresholds_1_address0;
reg    threshs_m_thresholds_1_ce0;
wire   [15:0] threshs_m_thresholds_1_q0;
wire   [3:0] threshs_m_thresholds_address0;
reg    threshs_m_thresholds_ce0;
wire   [15:0] threshs_m_thresholds_q0;
wire   [3:0] threshs_m_thresholds_11_address0;
reg    threshs_m_thresholds_11_ce0;
wire   [15:0] threshs_m_thresholds_11_q0;
wire   [3:0] threshs_m_thresholds_10_address0;
reg    threshs_m_thresholds_10_ce0;
wire   [15:0] threshs_m_thresholds_10_q0;
wire   [3:0] threshs_m_thresholds_9_address0;
reg    threshs_m_thresholds_9_ce0;
wire   [15:0] threshs_m_thresholds_9_q0;
wire   [3:0] threshs_m_thresholds_8_address0;
reg    threshs_m_thresholds_8_ce0;
wire   [15:0] threshs_m_thresholds_8_q0;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln248_fu_1079_p2;
wire   [0:0] icmp_ln252_fu_1094_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter3;
reg   [0:0] icmp_ln289_reg_3519;
reg   [0:0] icmp_ln289_reg_3519_pp0_iter2_reg;
reg    weight_V_V_TDATA_blk_n;
reg   [16:0] i_0_reg_1049;
reg    ap_predicate_op51_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
reg    ap_block_state5_io;
reg    ap_block_pp0_stage0_11001;
wire   [16:0] i_fu_1085_p2;
wire   [23:0] inElem_V_fu_1134_p11;
wire   [0:0] icmp_ln271_fu_1468_p2;
reg   [0:0] icmp_ln271_reg_3451;
reg   [0:0] icmp_ln271_reg_3451_pp0_iter1_reg;
wire   [3:0] trunc_ln647_fu_1474_p1;
reg  signed [3:0] trunc_ln647_reg_3459;
reg  signed [3:0] p_Result_1_0_1_reg_3464;
reg  signed [3:0] p_Result_1_0_2_reg_3469;
reg  signed [3:0] p_Result_1_1_reg_3474;
reg  signed [3:0] p_Result_1_1_1_reg_3479;
reg  signed [3:0] p_Result_1_1_2_reg_3484;
reg  signed [3:0] p_Result_1_2_reg_3489;
reg  signed [3:0] p_Result_1_2_1_reg_3494;
reg  signed [3:0] p_Result_1_2_2_reg_3499;
reg  signed [3:0] p_Result_1_3_reg_3504;
reg  signed [3:0] p_Result_1_3_1_reg_3509;
reg  signed [3:0] p_Result_1_3_2_reg_3514;
wire   [0:0] icmp_ln289_fu_1594_p2;
reg   [0:0] icmp_ln289_reg_3519_pp0_iter1_reg;
wire  signed [11:0] mul_ln1352_fu_1616_p2;
reg  signed [11:0] mul_ln1352_reg_3523;
wire   [12:0] add_ln700_1_fu_1676_p2;
reg   [12:0] add_ln700_1_reg_3528;
wire  signed [11:0] mul_ln1352_3_fu_1685_p2;
reg  signed [11:0] mul_ln1352_3_reg_3533;
wire   [12:0] add_ln700_4_fu_1717_p2;
reg   [12:0] add_ln700_4_reg_3538;
wire  signed [11:0] mul_ln1352_6_fu_1726_p2;
reg  signed [11:0] mul_ln1352_6_reg_3543;
wire   [12:0] add_ln700_7_fu_1758_p2;
reg   [12:0] add_ln700_7_reg_3548;
wire  signed [11:0] mul_ln1352_9_fu_1767_p2;
reg  signed [11:0] mul_ln1352_9_reg_3553;
wire   [12:0] add_ln700_10_fu_1799_p2;
reg   [12:0] add_ln700_10_reg_3558;
wire   [0:0] icmp_ln899_fu_2025_p2;
reg   [0:0] icmp_ln899_reg_3843;
wire   [0:0] icmp_ln899_1_fu_2031_p2;
reg   [0:0] icmp_ln899_1_reg_3848;
wire   [0:0] icmp_ln899_2_fu_2037_p2;
reg   [0:0] icmp_ln899_2_reg_3853;
wire   [0:0] icmp_ln899_3_fu_2043_p2;
reg   [0:0] icmp_ln899_3_reg_3858;
wire   [0:0] icmp_ln899_4_fu_2049_p2;
reg   [0:0] icmp_ln899_4_reg_3863;
wire   [0:0] icmp_ln899_5_fu_2055_p2;
reg   [0:0] icmp_ln899_5_reg_3868;
wire   [0:0] icmp_ln899_6_fu_2061_p2;
reg   [0:0] icmp_ln899_6_reg_3873;
wire   [0:0] xor_ln899_7_fu_2073_p2;
reg   [0:0] xor_ln899_7_reg_3878;
wire   [0:0] xor_ln899_8_fu_2085_p2;
reg   [0:0] xor_ln899_8_reg_3883;
wire   [0:0] xor_ln899_9_fu_2097_p2;
reg   [0:0] xor_ln899_9_reg_3888;
wire   [0:0] icmp_ln899_10_fu_2103_p2;
reg   [0:0] icmp_ln899_10_reg_3893;
wire   [0:0] icmp_ln899_11_fu_2109_p2;
reg   [0:0] icmp_ln899_11_reg_3898;
wire   [0:0] icmp_ln899_12_fu_2115_p2;
reg   [0:0] icmp_ln899_12_reg_3903;
wire   [0:0] icmp_ln899_13_fu_2121_p2;
reg   [0:0] icmp_ln899_13_reg_3908;
wire   [0:0] icmp_ln899_14_fu_2127_p2;
reg   [0:0] icmp_ln899_14_reg_3913;
wire   [0:0] icmp_ln899_15_fu_2133_p2;
reg   [0:0] icmp_ln899_15_reg_3918;
wire   [0:0] icmp_ln899_16_fu_2139_p2;
reg   [0:0] icmp_ln899_16_reg_3923;
wire   [0:0] icmp_ln899_17_fu_2145_p2;
reg   [0:0] icmp_ln899_17_reg_3928;
wire   [0:0] icmp_ln899_18_fu_2151_p2;
reg   [0:0] icmp_ln899_18_reg_3933;
wire   [0:0] icmp_ln899_19_fu_2157_p2;
reg   [0:0] icmp_ln899_19_reg_3938;
wire   [0:0] icmp_ln899_20_fu_2163_p2;
reg   [0:0] icmp_ln899_20_reg_3943;
wire   [0:0] xor_ln899_21_fu_2175_p2;
reg   [0:0] xor_ln899_21_reg_3948;
wire   [0:0] xor_ln899_22_fu_2187_p2;
reg   [0:0] xor_ln899_22_reg_3953;
wire   [0:0] xor_ln899_23_fu_2199_p2;
reg   [0:0] xor_ln899_23_reg_3958;
wire   [0:0] icmp_ln899_24_fu_2205_p2;
reg   [0:0] icmp_ln899_24_reg_3963;
wire   [0:0] icmp_ln899_25_fu_2211_p2;
reg   [0:0] icmp_ln899_25_reg_3968;
wire   [0:0] icmp_ln899_26_fu_2217_p2;
reg   [0:0] icmp_ln899_26_reg_3973;
wire   [0:0] icmp_ln899_27_fu_2223_p2;
reg   [0:0] icmp_ln899_27_reg_3978;
wire   [0:0] icmp_ln899_28_fu_2229_p2;
reg   [0:0] icmp_ln899_28_reg_3983;
wire   [0:0] icmp_ln899_29_fu_2235_p2;
reg   [0:0] icmp_ln899_29_reg_3988;
wire   [0:0] icmp_ln899_30_fu_2241_p2;
reg   [0:0] icmp_ln899_30_reg_3993;
wire   [0:0] icmp_ln899_31_fu_2247_p2;
reg   [0:0] icmp_ln899_31_reg_3998;
wire   [0:0] icmp_ln899_32_fu_2253_p2;
reg   [0:0] icmp_ln899_32_reg_4003;
wire   [0:0] icmp_ln899_33_fu_2259_p2;
reg   [0:0] icmp_ln899_33_reg_4008;
wire   [0:0] icmp_ln899_34_fu_2265_p2;
reg   [0:0] icmp_ln899_34_reg_4013;
wire   [0:0] xor_ln899_35_fu_2277_p2;
reg   [0:0] xor_ln899_35_reg_4018;
wire   [0:0] xor_ln899_36_fu_2289_p2;
reg   [0:0] xor_ln899_36_reg_4023;
wire   [0:0] xor_ln899_37_fu_2301_p2;
reg   [0:0] xor_ln899_37_reg_4028;
wire   [0:0] icmp_ln899_38_fu_2307_p2;
reg   [0:0] icmp_ln899_38_reg_4033;
wire   [0:0] icmp_ln899_39_fu_2313_p2;
reg   [0:0] icmp_ln899_39_reg_4038;
wire   [0:0] icmp_ln899_40_fu_2319_p2;
reg   [0:0] icmp_ln899_40_reg_4043;
wire   [0:0] icmp_ln899_41_fu_2325_p2;
reg   [0:0] icmp_ln899_41_reg_4048;
wire   [0:0] icmp_ln899_42_fu_2331_p2;
reg   [0:0] icmp_ln899_42_reg_4053;
wire   [0:0] icmp_ln899_43_fu_2337_p2;
reg   [0:0] icmp_ln899_43_reg_4058;
wire   [0:0] icmp_ln899_44_fu_2343_p2;
reg   [0:0] icmp_ln899_44_reg_4063;
wire   [0:0] icmp_ln899_45_fu_2349_p2;
reg   [0:0] icmp_ln899_45_reg_4068;
wire   [0:0] icmp_ln899_46_fu_2355_p2;
reg   [0:0] icmp_ln899_46_reg_4073;
wire   [0:0] icmp_ln899_47_fu_2361_p2;
reg   [0:0] icmp_ln899_47_reg_4078;
wire   [0:0] icmp_ln899_48_fu_2367_p2;
reg   [0:0] icmp_ln899_48_reg_4083;
wire   [0:0] xor_ln899_49_fu_2379_p2;
reg   [0:0] xor_ln899_49_reg_4088;
wire   [0:0] xor_ln899_50_fu_2391_p2;
reg   [0:0] xor_ln899_50_reg_4093;
wire   [0:0] xor_ln899_51_fu_2403_p2;
reg   [0:0] xor_ln899_51_reg_4098;
wire   [0:0] icmp_ln899_52_fu_2409_p2;
reg   [0:0] icmp_ln899_52_reg_4103;
wire   [0:0] icmp_ln899_53_fu_2415_p2;
reg   [0:0] icmp_ln899_53_reg_4108;
wire   [0:0] icmp_ln899_54_fu_2421_p2;
reg   [0:0] icmp_ln899_54_reg_4113;
wire   [0:0] icmp_ln899_55_fu_2427_p2;
reg   [0:0] icmp_ln899_55_reg_4118;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
wire   [23:0] ap_phi_reg_pp0_iter0_act_m_val_V_reg_1060;
reg   [23:0] ap_phi_reg_pp0_iter1_act_m_val_V_reg_1060;
wire   [63:0] zext_ln142_fu_1808_p1;
reg   [15:0] accu_V_0_0_0_fu_242;
wire   [15:0] accu_0_0_V_fu_1945_p2;
reg   [15:0] accu_V_0_1_0_fu_246;
wire   [15:0] accu_0_1_V_fu_1963_p2;
reg   [15:0] accu_V_0_2_0_fu_250;
wire   [15:0] accu_0_2_V_fu_1981_p2;
reg   [15:0] accu_V_0_3_0_fu_254;
wire   [15:0] accu_0_3_V_fu_1999_p2;
reg   [31:0] sf_1_fu_258;
wire   [31:0] sf_fu_1588_p2;
reg   [31:0] nf_assign_fu_262;
wire   [31:0] select_ln301_fu_1880_p3;
reg   [31:0] ap_sig_allocacmp_nf_assign_load_1;
reg   [23:0] inputBuf_8_V_1_fu_266;
wire   [23:0] inputBuf_8_V_19_fu_1412_p3;
reg   [23:0] inputBuf_8_V_2_fu_270;
wire   [23:0] inputBuf_8_V_18_fu_1404_p3;
reg   [23:0] inputBuf_8_V_4_fu_274;
wire   [23:0] inputBuf_8_V_16_fu_1388_p3;
reg   [23:0] inputBuf_8_V_6_fu_278;
wire   [23:0] inputBuf_8_V_15_fu_1372_p3;
reg   [23:0] inputBuf_8_V_7_fu_282;
wire   [23:0] inputBuf_8_V_14_fu_1348_p3;
reg   [23:0] inputBuf_8_V_5_fu_286;
wire   [23:0] inputBuf_8_V_13_fu_1332_p3;
reg   [23:0] inputBuf_8_V_3_fu_290;
wire   [23:0] inputBuf_8_V_12_fu_1308_p3;
reg   [23:0] inputBuf_8_V_8_fu_294;
wire   [23:0] inputBuf_8_V_11_fu_1284_p3;
reg   [23:0] inputBuf_8_V_9_fu_298;
wire   [23:0] inputBuf_8_V_fu_1252_p3;
reg    ap_block_pp0_stage0_01001;
wire   [3:0] inElem_V_fu_1134_p10;
wire   [3:0] trunc_ln321_fu_1158_p1;
wire   [0:0] icmp_ln321_7_fu_1204_p2;
wire   [0:0] icmp_ln321_6_fu_1198_p2;
wire   [0:0] icmp_ln321_5_fu_1192_p2;
wire   [0:0] icmp_ln321_4_fu_1186_p2;
wire   [0:0] icmp_ln321_3_fu_1180_p2;
wire   [0:0] icmp_ln321_2_fu_1174_p2;
wire   [0:0] icmp_ln321_1_fu_1168_p2;
wire   [0:0] icmp_ln321_fu_1162_p2;
wire   [0:0] or_ln321_fu_1210_p2;
wire   [0:0] or_ln321_1_fu_1216_p2;
wire   [0:0] or_ln321_2_fu_1222_p2;
wire   [0:0] or_ln321_3_fu_1228_p2;
wire   [0:0] or_ln321_4_fu_1234_p2;
wire   [0:0] or_ln321_5_fu_1240_p2;
wire   [0:0] or_ln321_6_fu_1246_p2;
wire   [23:0] select_ln321_fu_1260_p3;
wire   [23:0] select_ln321_1_fu_1268_p3;
wire   [23:0] select_ln321_2_fu_1276_p3;
wire   [23:0] select_ln321_4_fu_1292_p3;
wire   [23:0] select_ln321_5_fu_1300_p3;
wire   [23:0] select_ln321_7_fu_1316_p3;
wire   [23:0] select_ln321_8_fu_1324_p3;
wire   [23:0] select_ln321_10_fu_1340_p3;
wire   [23:0] select_ln321_12_fu_1356_p3;
wire   [23:0] select_ln321_13_fu_1364_p3;
wire   [23:0] select_ln321_15_fu_1380_p3;
wire   [23:0] inputBuf_8_V_17_fu_1396_p3;
wire   [7:0] trunc_ln647_1_fu_1605_p1;
wire  signed [7:0] mul_ln1352_fu_1616_p0;
wire  signed [11:0] sext_ln215_1_fu_1612_p1;
wire   [7:0] arg_V_read_assign_1_fu_1622_p4;
wire  signed [7:0] mul_ln1352_1_fu_1639_p0;
wire  signed [11:0] sext_ln215_3_fu_1635_p1;
wire  signed [11:0] mul_ln1352_1_fu_1639_p2;
wire   [7:0] arg_V_read_assign_2_fu_1649_p4;
wire  signed [7:0] mul_ln1352_2_fu_1666_p0;
wire  signed [11:0] sext_ln215_5_fu_1662_p1;
wire  signed [11:0] mul_ln1352_2_fu_1666_p2;
wire  signed [12:0] sext_ln700_1_fu_1672_p1;
wire  signed [12:0] sext_ln170_fu_1645_p1;
wire  signed [7:0] mul_ln1352_3_fu_1685_p0;
wire  signed [7:0] mul_ln1352_4_fu_1694_p0;
wire  signed [11:0] mul_ln1352_4_fu_1694_p2;
wire  signed [7:0] mul_ln1352_5_fu_1707_p0;
wire  signed [11:0] mul_ln1352_5_fu_1707_p2;
wire  signed [12:0] sext_ln700_4_fu_1713_p1;
wire  signed [12:0] sext_ln170_1_fu_1700_p1;
wire  signed [7:0] mul_ln1352_6_fu_1726_p0;
wire  signed [7:0] mul_ln1352_7_fu_1735_p0;
wire  signed [11:0] mul_ln1352_7_fu_1735_p2;
wire  signed [7:0] mul_ln1352_8_fu_1748_p0;
wire  signed [11:0] mul_ln1352_8_fu_1748_p2;
wire  signed [12:0] sext_ln700_7_fu_1754_p1;
wire  signed [12:0] sext_ln170_2_fu_1741_p1;
wire  signed [7:0] mul_ln1352_9_fu_1767_p0;
wire  signed [7:0] mul_ln1352_10_fu_1776_p0;
wire  signed [11:0] mul_ln1352_10_fu_1776_p2;
wire  signed [7:0] mul_ln1352_11_fu_1789_p0;
wire  signed [11:0] mul_ln1352_11_fu_1789_p2;
wire  signed [12:0] sext_ln700_10_fu_1795_p1;
wire  signed [12:0] sext_ln170_3_fu_1782_p1;
wire   [31:0] nf_fu_1868_p2;
wire   [0:0] icmp_ln301_fu_1874_p2;
wire  signed [15:0] sext_ln700_fu_1933_p1;
wire   [15:0] select_ln271_3_fu_1926_p3;
wire   [15:0] add_ln700_fu_1936_p2;
wire  signed [15:0] sext_ln700_2_fu_1942_p1;
wire  signed [15:0] sext_ln700_3_fu_1951_p1;
wire   [15:0] select_ln271_2_fu_1919_p3;
wire   [15:0] add_ln700_3_fu_1954_p2;
wire  signed [15:0] sext_ln700_5_fu_1960_p1;
wire  signed [15:0] sext_ln700_6_fu_1969_p1;
wire   [15:0] select_ln271_1_fu_1912_p3;
wire   [15:0] add_ln700_6_fu_1972_p2;
wire  signed [15:0] sext_ln700_8_fu_1978_p1;
wire  signed [15:0] sext_ln700_9_fu_1987_p1;
wire   [15:0] select_ln271_fu_1905_p3;
wire   [15:0] add_ln700_9_fu_1990_p2;
wire  signed [15:0] sext_ln700_11_fu_1996_p1;
wire   [0:0] icmp_ln899_7_fu_2067_p2;
wire   [0:0] icmp_ln899_8_fu_2079_p2;
wire   [0:0] icmp_ln899_9_fu_2091_p2;
wire   [0:0] icmp_ln899_21_fu_2169_p2;
wire   [0:0] icmp_ln899_22_fu_2181_p2;
wire   [0:0] icmp_ln899_23_fu_2193_p2;
wire   [0:0] icmp_ln899_35_fu_2271_p2;
wire   [0:0] icmp_ln899_36_fu_2283_p2;
wire   [0:0] icmp_ln899_37_fu_2295_p2;
wire   [0:0] icmp_ln899_49_fu_2373_p2;
wire   [0:0] icmp_ln899_50_fu_2385_p2;
wire   [0:0] icmp_ln899_51_fu_2397_p2;
wire   [0:0] xor_ln899_fu_2433_p2;
wire   [0:0] xor_ln899_1_fu_2446_p2;
wire   [0:0] xor_ln899_2_fu_2455_p2;
wire   [0:0] xor_ln899_3_fu_2464_p2;
wire   [0:0] xor_ln899_4_fu_2473_p2;
wire   [0:0] xor_ln899_5_fu_2482_p2;
wire   [0:0] xor_ln899_6_fu_2491_p2;
wire   [0:0] xor_ln899_10_fu_2509_p2;
wire   [0:0] xor_ln899_11_fu_2518_p2;
wire   [0:0] xor_ln899_12_fu_2527_p2;
wire   [0:0] xor_ln899_13_fu_2536_p2;
wire   [1:0] zext_ln142_1_fu_2451_p1;
wire   [1:0] zext_ln142_2_fu_2460_p1;
wire   [1:0] add_ln700_12_fu_2545_p2;
wire   [3:0] zext_ln700_1_fu_2551_p1;
wire   [3:0] select_ln700_fu_2438_p3;
wire   [1:0] zext_ln142_3_fu_2469_p1;
wire   [1:0] zext_ln142_4_fu_2478_p1;
wire   [1:0] add_ln700_14_fu_2561_p2;
wire   [1:0] zext_ln142_5_fu_2487_p1;
wire   [1:0] zext_ln142_6_fu_2496_p1;
wire   [1:0] add_ln700_15_fu_2571_p2;
wire   [2:0] zext_ln700_3_fu_2577_p1;
wire   [2:0] zext_ln700_2_fu_2567_p1;
wire   [2:0] add_ln700_16_fu_2581_p2;
wire   [3:0] zext_ln700_4_fu_2587_p1;
wire   [3:0] add_ln700_13_fu_2555_p2;
wire   [1:0] zext_ln142_8_fu_2503_p1;
wire   [1:0] zext_ln142_9_fu_2506_p1;
wire   [1:0] add_ln700_18_fu_2597_p2;
wire   [1:0] zext_ln142_7_fu_2500_p1;
wire   [1:0] add_ln700_19_fu_2603_p2;
wire   [1:0] zext_ln142_10_fu_2514_p1;
wire   [1:0] zext_ln142_11_fu_2523_p1;
wire   [1:0] add_ln700_20_fu_2613_p2;
wire   [1:0] zext_ln142_12_fu_2532_p1;
wire   [1:0] zext_ln700_fu_2541_p1;
wire   [1:0] add_ln700_21_fu_2623_p2;
wire   [2:0] zext_ln700_7_fu_2629_p1;
wire   [2:0] zext_ln700_6_fu_2619_p1;
wire   [2:0] add_ln700_22_fu_2633_p2;
wire   [2:0] zext_ln700_5_fu_2609_p1;
wire   [2:0] add_ln700_23_fu_2639_p2;
wire   [3:0] zext_ln700_8_fu_2645_p1;
wire   [3:0] add_ln700_17_fu_2591_p2;
wire   [0:0] xor_ln899_14_fu_2655_p2;
wire   [0:0] xor_ln899_15_fu_2668_p2;
wire   [0:0] xor_ln899_16_fu_2677_p2;
wire   [0:0] xor_ln899_17_fu_2686_p2;
wire   [0:0] xor_ln899_18_fu_2695_p2;
wire   [0:0] xor_ln899_19_fu_2704_p2;
wire   [0:0] xor_ln899_20_fu_2713_p2;
wire   [0:0] xor_ln899_24_fu_2731_p2;
wire   [0:0] xor_ln899_25_fu_2740_p2;
wire   [0:0] xor_ln899_26_fu_2749_p2;
wire   [0:0] xor_ln899_27_fu_2758_p2;
wire   [1:0] zext_ln142_13_fu_2673_p1;
wire   [1:0] zext_ln142_14_fu_2682_p1;
wire   [1:0] add_ln700_25_fu_2767_p2;
wire   [3:0] zext_ln700_10_fu_2773_p1;
wire   [3:0] select_ln700_1_fu_2660_p3;
wire   [1:0] zext_ln142_15_fu_2691_p1;
wire   [1:0] zext_ln142_16_fu_2700_p1;
wire   [1:0] add_ln700_27_fu_2783_p2;
wire   [1:0] zext_ln142_17_fu_2709_p1;
wire   [1:0] zext_ln142_18_fu_2718_p1;
wire   [1:0] add_ln700_28_fu_2793_p2;
wire   [2:0] zext_ln700_12_fu_2799_p1;
wire   [2:0] zext_ln700_11_fu_2789_p1;
wire   [2:0] add_ln700_29_fu_2803_p2;
wire   [3:0] zext_ln700_13_fu_2809_p1;
wire   [3:0] add_ln700_26_fu_2777_p2;
wire   [1:0] zext_ln142_20_fu_2725_p1;
wire   [1:0] zext_ln142_21_fu_2728_p1;
wire   [1:0] add_ln700_31_fu_2819_p2;
wire   [1:0] zext_ln142_19_fu_2722_p1;
wire   [1:0] add_ln700_32_fu_2825_p2;
wire   [1:0] zext_ln142_22_fu_2736_p1;
wire   [1:0] zext_ln142_23_fu_2745_p1;
wire   [1:0] add_ln700_33_fu_2835_p2;
wire   [1:0] zext_ln142_24_fu_2754_p1;
wire   [1:0] zext_ln700_9_fu_2763_p1;
wire   [1:0] add_ln700_34_fu_2845_p2;
wire   [2:0] zext_ln700_16_fu_2851_p1;
wire   [2:0] zext_ln700_15_fu_2841_p1;
wire   [2:0] add_ln700_35_fu_2855_p2;
wire   [2:0] zext_ln700_14_fu_2831_p1;
wire   [2:0] add_ln700_36_fu_2861_p2;
wire   [3:0] zext_ln700_17_fu_2867_p1;
wire   [3:0] add_ln700_30_fu_2813_p2;
wire   [0:0] xor_ln899_28_fu_2877_p2;
wire   [0:0] xor_ln899_29_fu_2890_p2;
wire   [0:0] xor_ln899_30_fu_2899_p2;
wire   [0:0] xor_ln899_31_fu_2908_p2;
wire   [0:0] xor_ln899_32_fu_2917_p2;
wire   [0:0] xor_ln899_33_fu_2926_p2;
wire   [0:0] xor_ln899_34_fu_2935_p2;
wire   [0:0] xor_ln899_38_fu_2953_p2;
wire   [0:0] xor_ln899_39_fu_2962_p2;
wire   [0:0] xor_ln899_40_fu_2971_p2;
wire   [0:0] xor_ln899_41_fu_2980_p2;
wire   [1:0] zext_ln142_25_fu_2895_p1;
wire   [1:0] zext_ln142_26_fu_2904_p1;
wire   [1:0] add_ln700_38_fu_2989_p2;
wire   [3:0] zext_ln700_19_fu_2995_p1;
wire   [3:0] select_ln700_2_fu_2882_p3;
wire   [1:0] zext_ln142_27_fu_2913_p1;
wire   [1:0] zext_ln142_28_fu_2922_p1;
wire   [1:0] add_ln700_40_fu_3005_p2;
wire   [1:0] zext_ln142_29_fu_2931_p1;
wire   [1:0] zext_ln142_30_fu_2940_p1;
wire   [1:0] add_ln700_41_fu_3015_p2;
wire   [2:0] zext_ln700_21_fu_3021_p1;
wire   [2:0] zext_ln700_20_fu_3011_p1;
wire   [2:0] add_ln700_42_fu_3025_p2;
wire   [3:0] zext_ln700_22_fu_3031_p1;
wire   [3:0] add_ln700_39_fu_2999_p2;
wire   [1:0] zext_ln142_32_fu_2947_p1;
wire   [1:0] zext_ln142_33_fu_2950_p1;
wire   [1:0] add_ln700_44_fu_3041_p2;
wire   [1:0] zext_ln142_31_fu_2944_p1;
wire   [1:0] add_ln700_45_fu_3047_p2;
wire   [1:0] zext_ln142_34_fu_2958_p1;
wire   [1:0] zext_ln142_35_fu_2967_p1;
wire   [1:0] add_ln700_46_fu_3057_p2;
wire   [1:0] zext_ln142_36_fu_2976_p1;
wire   [1:0] zext_ln700_18_fu_2985_p1;
wire   [1:0] add_ln700_47_fu_3067_p2;
wire   [2:0] zext_ln700_25_fu_3073_p1;
wire   [2:0] zext_ln700_24_fu_3063_p1;
wire   [2:0] add_ln700_48_fu_3077_p2;
wire   [2:0] zext_ln700_23_fu_3053_p1;
wire   [2:0] add_ln700_49_fu_3083_p2;
wire   [3:0] zext_ln700_26_fu_3089_p1;
wire   [3:0] add_ln700_43_fu_3035_p2;
wire   [0:0] xor_ln899_42_fu_3099_p2;
wire   [0:0] xor_ln899_43_fu_3112_p2;
wire   [0:0] xor_ln899_44_fu_3121_p2;
wire   [0:0] xor_ln899_45_fu_3130_p2;
wire   [0:0] xor_ln899_46_fu_3139_p2;
wire   [0:0] xor_ln899_47_fu_3148_p2;
wire   [0:0] xor_ln899_48_fu_3157_p2;
wire   [0:0] xor_ln899_52_fu_3175_p2;
wire   [0:0] xor_ln899_53_fu_3184_p2;
wire   [0:0] xor_ln899_54_fu_3193_p2;
wire   [0:0] xor_ln899_55_fu_3202_p2;
wire   [1:0] zext_ln142_37_fu_3117_p1;
wire   [1:0] zext_ln142_38_fu_3126_p1;
wire   [1:0] add_ln700_51_fu_3211_p2;
wire   [3:0] zext_ln700_28_fu_3217_p1;
wire   [3:0] select_ln700_3_fu_3104_p3;
wire   [1:0] zext_ln142_39_fu_3135_p1;
wire   [1:0] zext_ln142_40_fu_3144_p1;
wire   [1:0] add_ln700_53_fu_3227_p2;
wire   [1:0] zext_ln142_41_fu_3153_p1;
wire   [1:0] zext_ln142_42_fu_3162_p1;
wire   [1:0] add_ln700_54_fu_3237_p2;
wire   [2:0] zext_ln700_30_fu_3243_p1;
wire   [2:0] zext_ln700_29_fu_3233_p1;
wire   [2:0] add_ln700_55_fu_3247_p2;
wire   [3:0] zext_ln700_31_fu_3253_p1;
wire   [3:0] add_ln700_52_fu_3221_p2;
wire   [1:0] zext_ln142_44_fu_3169_p1;
wire   [1:0] zext_ln142_45_fu_3172_p1;
wire   [1:0] add_ln700_57_fu_3263_p2;
wire   [1:0] zext_ln142_43_fu_3166_p1;
wire   [1:0] add_ln700_58_fu_3269_p2;
wire   [1:0] zext_ln142_46_fu_3180_p1;
wire   [1:0] zext_ln142_47_fu_3189_p1;
wire   [1:0] add_ln700_59_fu_3279_p2;
wire   [1:0] zext_ln142_48_fu_3198_p1;
wire   [1:0] zext_ln700_27_fu_3207_p1;
wire   [1:0] add_ln700_60_fu_3289_p2;
wire   [2:0] zext_ln700_34_fu_3295_p1;
wire   [2:0] zext_ln700_33_fu_3285_p1;
wire   [2:0] add_ln700_61_fu_3299_p2;
wire   [2:0] zext_ln700_32_fu_3275_p1;
wire   [2:0] add_ln700_62_fu_3305_p2;
wire   [3:0] zext_ln700_35_fu_3311_p1;
wire   [3:0] add_ln700_56_fu_3257_p2;
wire   [3:0] add_ln700_63_fu_3315_p2;
wire   [3:0] add_ln700_50_fu_3093_p2;
wire   [3:0] add_ln700_37_fu_2871_p2;
wire   [3:0] add_ln700_24_fu_2649_p2;
wire    ap_CS_fsm_state6;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_485;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

StreamingFCLayer_Batch_2_Matrix_Vector_Actbkb #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_55_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_55_address0),
    .ce0(threshs_m_thresholds_55_ce0),
    .q0(threshs_m_thresholds_55_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actcud #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_54_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_54_address0),
    .ce0(threshs_m_thresholds_54_ce0),
    .q0(threshs_m_thresholds_54_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActdEe #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_49_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_49_address0),
    .ce0(threshs_m_thresholds_49_ce0),
    .q0(threshs_m_thresholds_49_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActeOg #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_48_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_48_address0),
    .ce0(threshs_m_thresholds_48_ce0),
    .q0(threshs_m_thresholds_48_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActfYi #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_47_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_47_address0),
    .ce0(threshs_m_thresholds_47_ce0),
    .q0(threshs_m_thresholds_47_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actg8j #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_46_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_46_address0),
    .ce0(threshs_m_thresholds_46_ce0),
    .q0(threshs_m_thresholds_46_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Acthbi #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_45_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_45_address0),
    .ce0(threshs_m_thresholds_45_ce0),
    .q0(threshs_m_thresholds_45_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actibs #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_44_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_44_address0),
    .ce0(threshs_m_thresholds_44_ce0),
    .q0(threshs_m_thresholds_44_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActjbC #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_43_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_43_address0),
    .ce0(threshs_m_thresholds_43_ce0),
    .q0(threshs_m_thresholds_43_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActkbM #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_42_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_42_address0),
    .ce0(threshs_m_thresholds_42_ce0),
    .q0(threshs_m_thresholds_42_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActlbW #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_53_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_53_address0),
    .ce0(threshs_m_thresholds_53_ce0),
    .q0(threshs_m_thresholds_53_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actmb6 #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_52_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_52_address0),
    .ce0(threshs_m_thresholds_52_ce0),
    .q0(threshs_m_thresholds_52_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actncg #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_51_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_51_address0),
    .ce0(threshs_m_thresholds_51_ce0),
    .q0(threshs_m_thresholds_51_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actocq #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_50_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_50_address0),
    .ce0(threshs_m_thresholds_50_ce0),
    .q0(threshs_m_thresholds_50_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActpcA #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_41_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_41_address0),
    .ce0(threshs_m_thresholds_41_ce0),
    .q0(threshs_m_thresholds_41_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActqcK #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_40_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_40_address0),
    .ce0(threshs_m_thresholds_40_ce0),
    .q0(threshs_m_thresholds_40_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActrcU #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_35_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_35_address0),
    .ce0(threshs_m_thresholds_35_ce0),
    .q0(threshs_m_thresholds_35_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actsc4 #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_34_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_34_address0),
    .ce0(threshs_m_thresholds_34_ce0),
    .q0(threshs_m_thresholds_34_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Acttde #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_33_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_33_address0),
    .ce0(threshs_m_thresholds_33_ce0),
    .q0(threshs_m_thresholds_33_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actudo #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_32_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_32_address0),
    .ce0(threshs_m_thresholds_32_ce0),
    .q0(threshs_m_thresholds_32_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actvdy #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_31_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_31_address0),
    .ce0(threshs_m_thresholds_31_ce0),
    .q0(threshs_m_thresholds_31_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActwdI #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_30_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_30_address0),
    .ce0(threshs_m_thresholds_30_ce0),
    .q0(threshs_m_thresholds_30_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActxdS #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_29_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_29_address0),
    .ce0(threshs_m_thresholds_29_ce0),
    .q0(threshs_m_thresholds_29_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actyd2 #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_28_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_28_address0),
    .ce0(threshs_m_thresholds_28_ce0),
    .q0(threshs_m_thresholds_28_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Actzec #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_39_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_39_address0),
    .ce0(threshs_m_thresholds_39_ce0),
    .q0(threshs_m_thresholds_39_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActAem #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_38_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_38_address0),
    .ce0(threshs_m_thresholds_38_ce0),
    .q0(threshs_m_thresholds_38_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActBew #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_37_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_37_address0),
    .ce0(threshs_m_thresholds_37_ce0),
    .q0(threshs_m_thresholds_37_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActCeG #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_36_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_36_address0),
    .ce0(threshs_m_thresholds_36_ce0),
    .q0(threshs_m_thresholds_36_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActDeQ #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_27_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_27_address0),
    .ce0(threshs_m_thresholds_27_ce0),
    .q0(threshs_m_thresholds_27_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActEe0 #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_26_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_26_address0),
    .ce0(threshs_m_thresholds_26_ce0),
    .q0(threshs_m_thresholds_26_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActFfa #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_21_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_21_address0),
    .ce0(threshs_m_thresholds_21_ce0),
    .q0(threshs_m_thresholds_21_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActGfk #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_20_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_20_address0),
    .ce0(threshs_m_thresholds_20_ce0),
    .q0(threshs_m_thresholds_20_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActHfu #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_19_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_19_address0),
    .ce0(threshs_m_thresholds_19_ce0),
    .q0(threshs_m_thresholds_19_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActHfu #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_18_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_18_address0),
    .ce0(threshs_m_thresholds_18_ce0),
    .q0(threshs_m_thresholds_18_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActHfu #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_17_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_17_address0),
    .ce0(threshs_m_thresholds_17_ce0),
    .q0(threshs_m_thresholds_17_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActHfu #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_16_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_16_address0),
    .ce0(threshs_m_thresholds_16_ce0),
    .q0(threshs_m_thresholds_16_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActLf8 #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_15_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_15_address0),
    .ce0(threshs_m_thresholds_15_ce0),
    .q0(threshs_m_thresholds_15_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActMgi #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_14_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_14_address0),
    .ce0(threshs_m_thresholds_14_ce0),
    .q0(threshs_m_thresholds_14_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActNgs #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_25_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_25_address0),
    .ce0(threshs_m_thresholds_25_ce0),
    .q0(threshs_m_thresholds_25_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActOgC #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_24_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_24_address0),
    .ce0(threshs_m_thresholds_24_ce0),
    .q0(threshs_m_thresholds_24_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActPgM #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_23_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_23_address0),
    .ce0(threshs_m_thresholds_23_ce0),
    .q0(threshs_m_thresholds_23_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActQgW #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_22_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_22_address0),
    .ce0(threshs_m_thresholds_22_ce0),
    .q0(threshs_m_thresholds_22_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActRg6 #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_13_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_13_address0),
    .ce0(threshs_m_thresholds_13_ce0),
    .q0(threshs_m_thresholds_13_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActShg #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_12_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_12_address0),
    .ce0(threshs_m_thresholds_12_ce0),
    .q0(threshs_m_thresholds_12_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActThq #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_7_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_7_address0),
    .ce0(threshs_m_thresholds_7_ce0),
    .q0(threshs_m_thresholds_7_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActUhA #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_6_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_6_address0),
    .ce0(threshs_m_thresholds_6_ce0),
    .q0(threshs_m_thresholds_6_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActVhK #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_5_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_5_address0),
    .ce0(threshs_m_thresholds_5_ce0),
    .q0(threshs_m_thresholds_5_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActWhU #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_4_address0),
    .ce0(threshs_m_thresholds_4_ce0),
    .q0(threshs_m_thresholds_4_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActXh4 #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_3_address0),
    .ce0(threshs_m_thresholds_3_ce0),
    .q0(threshs_m_thresholds_3_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActYie #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_2_address0),
    .ce0(threshs_m_thresholds_2_ce0),
    .q0(threshs_m_thresholds_2_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_ActZio #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_1_address0),
    .ce0(threshs_m_thresholds_1_ce0),
    .q0(threshs_m_thresholds_1_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Act0iy #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_address0),
    .ce0(threshs_m_thresholds_ce0),
    .q0(threshs_m_thresholds_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Act1iI #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_11_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_11_address0),
    .ce0(threshs_m_thresholds_11_ce0),
    .q0(threshs_m_thresholds_11_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Act2iS #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_10_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_10_address0),
    .ce0(threshs_m_thresholds_10_ce0),
    .q0(threshs_m_thresholds_10_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Act3i2 #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_9_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_9_address0),
    .ce0(threshs_m_thresholds_9_ce0),
    .q0(threshs_m_thresholds_9_q0)
);

StreamingFCLayer_Batch_2_Matrix_Vector_Act4jc #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
threshs_m_thresholds_8_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_8_address0),
    .ce0(threshs_m_thresholds_8_ce0),
    .q0(threshs_m_thresholds_8_q0)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_5jm #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 24 ),
    .din1_WIDTH( 24 ),
    .din2_WIDTH( 24 ),
    .din3_WIDTH( 24 ),
    .din4_WIDTH( 24 ),
    .din5_WIDTH( 24 ),
    .din6_WIDTH( 24 ),
    .din7_WIDTH( 24 ),
    .din8_WIDTH( 24 ),
    .din9_WIDTH( 4 ),
    .dout_WIDTH( 24 ))
StreamingFCLayer_5jm_U1(
    .din0(inputBuf_8_V_1_fu_266),
    .din1(inputBuf_8_V_2_fu_270),
    .din2(inputBuf_8_V_4_fu_274),
    .din3(inputBuf_8_V_6_fu_278),
    .din4(inputBuf_8_V_7_fu_282),
    .din5(inputBuf_8_V_5_fu_286),
    .din6(inputBuf_8_V_3_fu_290),
    .din7(inputBuf_8_V_8_fu_294),
    .din8(inputBuf_8_V_9_fu_298),
    .din9(inElem_V_fu_1134_p10),
    .dout(inElem_V_fu_1134_p11)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U2(
    .din0(mul_ln1352_fu_1616_p0),
    .din1(trunc_ln647_reg_3459),
    .dout(mul_ln1352_fu_1616_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U3(
    .din0(mul_ln1352_1_fu_1639_p0),
    .din1(p_Result_1_0_1_reg_3464),
    .dout(mul_ln1352_1_fu_1639_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U4(
    .din0(mul_ln1352_2_fu_1666_p0),
    .din1(p_Result_1_0_2_reg_3469),
    .dout(mul_ln1352_2_fu_1666_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U5(
    .din0(mul_ln1352_3_fu_1685_p0),
    .din1(p_Result_1_1_reg_3474),
    .dout(mul_ln1352_3_fu_1685_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U6(
    .din0(mul_ln1352_4_fu_1694_p0),
    .din1(p_Result_1_1_1_reg_3479),
    .dout(mul_ln1352_4_fu_1694_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U7(
    .din0(mul_ln1352_5_fu_1707_p0),
    .din1(p_Result_1_1_2_reg_3484),
    .dout(mul_ln1352_5_fu_1707_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U8(
    .din0(mul_ln1352_6_fu_1726_p0),
    .din1(p_Result_1_2_reg_3489),
    .dout(mul_ln1352_6_fu_1726_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U9(
    .din0(mul_ln1352_7_fu_1735_p0),
    .din1(p_Result_1_2_1_reg_3494),
    .dout(mul_ln1352_7_fu_1735_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U10(
    .din0(mul_ln1352_8_fu_1748_p0),
    .din1(p_Result_1_2_2_reg_3499),
    .dout(mul_ln1352_8_fu_1748_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U11(
    .din0(mul_ln1352_9_fu_1767_p0),
    .din1(p_Result_1_3_reg_3504),
    .dout(mul_ln1352_9_fu_1767_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U12(
    .din0(mul_ln1352_10_fu_1776_p0),
    .din1(p_Result_1_3_1_reg_3509),
    .dout(mul_ln1352_10_fu_1776_p2)
);

StreamingFCLayer_Batch_2_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 12 ))
StreamingFCLayer_6jw_U13(
    .din0(mul_ln1352_11_fu_1789_p0),
    .din1(p_Result_1_3_2_reg_3514),
    .dout(mul_ln1352_11_fu_1789_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_condition_485)) begin
        if (((icmp_ln252_fu_1094_p2 == 1'd0) & (icmp_ln248_fu_1079_p2 == 1'd0))) begin
            ap_phi_reg_pp0_iter1_act_m_val_V_reg_1060 <= inElem_V_fu_1134_p11;
        end else if (((icmp_ln252_fu_1094_p2 == 1'd1) & (icmp_ln248_fu_1079_p2 == 1'd0))) begin
            ap_phi_reg_pp0_iter1_act_m_val_V_reg_1060 <= in_V_V_TDATA;
        end else if ((1'b1 == 1'b1)) begin
            ap_phi_reg_pp0_iter1_act_m_val_V_reg_1060 <= ap_phi_reg_pp0_iter0_act_m_val_V_reg_1060;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_1079_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_reg_1049 <= i_fu_1085_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_reg_1049 <= 17'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_3519 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        nf_assign_fu_262 <= select_ln301_fu_1880_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        nf_assign_fu_262 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_1594_p2 == 1'd0) & (icmp_ln248_fu_1079_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        sf_1_fu_258 <= sf_fu_1588_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_1594_p2 == 1'd1) & (icmp_ln248_fu_1079_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        sf_1_fu_258 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        accu_V_0_0_0_fu_242 <= accu_0_0_V_fu_1945_p2;
        accu_V_0_1_0_fu_246 <= accu_0_1_V_fu_1963_p2;
        accu_V_0_2_0_fu_250 <= accu_0_2_V_fu_1981_p2;
        accu_V_0_3_0_fu_254 <= accu_0_3_V_fu_1999_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln700_10_reg_3558 <= add_ln700_10_fu_1799_p2;
        add_ln700_1_reg_3528 <= add_ln700_1_fu_1676_p2;
        add_ln700_4_reg_3538 <= add_ln700_4_fu_1717_p2;
        add_ln700_7_reg_3548 <= add_ln700_7_fu_1758_p2;
        icmp_ln271_reg_3451_pp0_iter1_reg <= icmp_ln271_reg_3451;
        icmp_ln289_reg_3519_pp0_iter1_reg <= icmp_ln289_reg_3519;
        mul_ln1352_3_reg_3533 <= mul_ln1352_3_fu_1685_p2;
        mul_ln1352_6_reg_3543 <= mul_ln1352_6_fu_1726_p2;
        mul_ln1352_9_reg_3553 <= mul_ln1352_9_fu_1767_p2;
        mul_ln1352_reg_3523 <= mul_ln1352_fu_1616_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_1079_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln271_reg_3451 <= icmp_ln271_fu_1468_p2;
        icmp_ln289_reg_3519 <= icmp_ln289_fu_1594_p2;
        p_Result_1_0_1_reg_3464 <= {{weight_V_V_TDATA[7:4]}};
        p_Result_1_0_2_reg_3469 <= {{weight_V_V_TDATA[11:8]}};
        p_Result_1_1_1_reg_3479 <= {{weight_V_V_TDATA[19:16]}};
        p_Result_1_1_2_reg_3484 <= {{weight_V_V_TDATA[23:20]}};
        p_Result_1_1_reg_3474 <= {{weight_V_V_TDATA[15:12]}};
        p_Result_1_2_1_reg_3494 <= {{weight_V_V_TDATA[31:28]}};
        p_Result_1_2_2_reg_3499 <= {{weight_V_V_TDATA[35:32]}};
        p_Result_1_2_reg_3489 <= {{weight_V_V_TDATA[27:24]}};
        p_Result_1_3_1_reg_3509 <= {{weight_V_V_TDATA[43:40]}};
        p_Result_1_3_2_reg_3514 <= {{weight_V_V_TDATA[47:44]}};
        p_Result_1_3_reg_3504 <= {{weight_V_V_TDATA[39:36]}};
        trunc_ln647_reg_3459 <= trunc_ln647_fu_1474_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln289_reg_3519_pp0_iter2_reg <= icmp_ln289_reg_3519_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_3519_pp0_iter1_reg == 1'd1))) begin
        icmp_ln899_10_reg_3893 <= icmp_ln899_10_fu_2103_p2;
        icmp_ln899_11_reg_3898 <= icmp_ln899_11_fu_2109_p2;
        icmp_ln899_12_reg_3903 <= icmp_ln899_12_fu_2115_p2;
        icmp_ln899_13_reg_3908 <= icmp_ln899_13_fu_2121_p2;
        icmp_ln899_14_reg_3913 <= icmp_ln899_14_fu_2127_p2;
        icmp_ln899_15_reg_3918 <= icmp_ln899_15_fu_2133_p2;
        icmp_ln899_16_reg_3923 <= icmp_ln899_16_fu_2139_p2;
        icmp_ln899_17_reg_3928 <= icmp_ln899_17_fu_2145_p2;
        icmp_ln899_18_reg_3933 <= icmp_ln899_18_fu_2151_p2;
        icmp_ln899_19_reg_3938 <= icmp_ln899_19_fu_2157_p2;
        icmp_ln899_1_reg_3848 <= icmp_ln899_1_fu_2031_p2;
        icmp_ln899_20_reg_3943 <= icmp_ln899_20_fu_2163_p2;
        icmp_ln899_24_reg_3963 <= icmp_ln899_24_fu_2205_p2;
        icmp_ln899_25_reg_3968 <= icmp_ln899_25_fu_2211_p2;
        icmp_ln899_26_reg_3973 <= icmp_ln899_26_fu_2217_p2;
        icmp_ln899_27_reg_3978 <= icmp_ln899_27_fu_2223_p2;
        icmp_ln899_28_reg_3983 <= icmp_ln899_28_fu_2229_p2;
        icmp_ln899_29_reg_3988 <= icmp_ln899_29_fu_2235_p2;
        icmp_ln899_2_reg_3853 <= icmp_ln899_2_fu_2037_p2;
        icmp_ln899_30_reg_3993 <= icmp_ln899_30_fu_2241_p2;
        icmp_ln899_31_reg_3998 <= icmp_ln899_31_fu_2247_p2;
        icmp_ln899_32_reg_4003 <= icmp_ln899_32_fu_2253_p2;
        icmp_ln899_33_reg_4008 <= icmp_ln899_33_fu_2259_p2;
        icmp_ln899_34_reg_4013 <= icmp_ln899_34_fu_2265_p2;
        icmp_ln899_38_reg_4033 <= icmp_ln899_38_fu_2307_p2;
        icmp_ln899_39_reg_4038 <= icmp_ln899_39_fu_2313_p2;
        icmp_ln899_3_reg_3858 <= icmp_ln899_3_fu_2043_p2;
        icmp_ln899_40_reg_4043 <= icmp_ln899_40_fu_2319_p2;
        icmp_ln899_41_reg_4048 <= icmp_ln899_41_fu_2325_p2;
        icmp_ln899_42_reg_4053 <= icmp_ln899_42_fu_2331_p2;
        icmp_ln899_43_reg_4058 <= icmp_ln899_43_fu_2337_p2;
        icmp_ln899_44_reg_4063 <= icmp_ln899_44_fu_2343_p2;
        icmp_ln899_45_reg_4068 <= icmp_ln899_45_fu_2349_p2;
        icmp_ln899_46_reg_4073 <= icmp_ln899_46_fu_2355_p2;
        icmp_ln899_47_reg_4078 <= icmp_ln899_47_fu_2361_p2;
        icmp_ln899_48_reg_4083 <= icmp_ln899_48_fu_2367_p2;
        icmp_ln899_4_reg_3863 <= icmp_ln899_4_fu_2049_p2;
        icmp_ln899_52_reg_4103 <= icmp_ln899_52_fu_2409_p2;
        icmp_ln899_53_reg_4108 <= icmp_ln899_53_fu_2415_p2;
        icmp_ln899_54_reg_4113 <= icmp_ln899_54_fu_2421_p2;
        icmp_ln899_55_reg_4118 <= icmp_ln899_55_fu_2427_p2;
        icmp_ln899_5_reg_3868 <= icmp_ln899_5_fu_2055_p2;
        icmp_ln899_6_reg_3873 <= icmp_ln899_6_fu_2061_p2;
        icmp_ln899_reg_3843 <= icmp_ln899_fu_2025_p2;
        xor_ln899_21_reg_3948 <= xor_ln899_21_fu_2175_p2;
        xor_ln899_22_reg_3953 <= xor_ln899_22_fu_2187_p2;
        xor_ln899_23_reg_3958 <= xor_ln899_23_fu_2199_p2;
        xor_ln899_35_reg_4018 <= xor_ln899_35_fu_2277_p2;
        xor_ln899_36_reg_4023 <= xor_ln899_36_fu_2289_p2;
        xor_ln899_37_reg_4028 <= xor_ln899_37_fu_2301_p2;
        xor_ln899_49_reg_4088 <= xor_ln899_49_fu_2379_p2;
        xor_ln899_50_reg_4093 <= xor_ln899_50_fu_2391_p2;
        xor_ln899_51_reg_4098 <= xor_ln899_51_fu_2403_p2;
        xor_ln899_7_reg_3878 <= xor_ln899_7_fu_2073_p2;
        xor_ln899_8_reg_3883 <= xor_ln899_8_fu_2085_p2;
        xor_ln899_9_reg_3888 <= xor_ln899_9_fu_2097_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1094_p2 == 1'd1) & (icmp_ln248_fu_1079_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_8_V_1_fu_266 <= inputBuf_8_V_19_fu_1412_p3;
        inputBuf_8_V_2_fu_270 <= inputBuf_8_V_18_fu_1404_p3;
        inputBuf_8_V_3_fu_290 <= inputBuf_8_V_12_fu_1308_p3;
        inputBuf_8_V_4_fu_274 <= inputBuf_8_V_16_fu_1388_p3;
        inputBuf_8_V_5_fu_286 <= inputBuf_8_V_13_fu_1332_p3;
        inputBuf_8_V_6_fu_278 <= inputBuf_8_V_15_fu_1372_p3;
        inputBuf_8_V_7_fu_282 <= inputBuf_8_V_14_fu_1348_p3;
        inputBuf_8_V_8_fu_294 <= inputBuf_8_V_11_fu_1284_p3;
        inputBuf_8_V_9_fu_298 <= inputBuf_8_V_fu_1252_p3;
    end
end

always @ (*) begin
    if ((icmp_ln248_fu_1079_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state6) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_3519 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_sig_allocacmp_nf_assign_load_1 = select_ln301_fu_1880_p3;
    end else begin
        ap_sig_allocacmp_nf_assign_load_1 = nf_assign_fu_262;
    end
end

always @ (*) begin
    if (((icmp_ln252_fu_1094_p2 == 1'd1) & (icmp_ln248_fu_1079_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op51_read_state2 == 1'b1))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_3519_pp0_iter2_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_3519_pp0_iter2_reg == 1'd1) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_10_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_10_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_11_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_11_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_12_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_12_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_13_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_13_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_14_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_14_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_15_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_15_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_16_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_16_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_17_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_17_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_18_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_18_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_19_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_19_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_1_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_1_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_20_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_20_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_21_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_21_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_22_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_22_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_23_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_23_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_24_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_24_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_25_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_25_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_26_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_26_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_27_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_27_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_28_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_28_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_29_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_29_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_2_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_2_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_30_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_30_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_31_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_31_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_32_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_32_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_33_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_33_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_34_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_34_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_35_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_35_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_36_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_36_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_37_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_37_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_38_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_38_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_39_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_39_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_3_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_3_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_40_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_40_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_41_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_41_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_42_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_42_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_43_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_43_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_44_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_44_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_45_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_45_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_46_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_46_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_47_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_47_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_48_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_48_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_49_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_49_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_4_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_4_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_50_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_50_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_51_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_51_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_52_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_52_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_53_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_53_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_54_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_54_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_55_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_55_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_5_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_5_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_6_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_6_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_7_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_7_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_8_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_8_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_9_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_9_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln248_fu_1079_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TDATA_blk_n = weight_V_V_TVALID;
    end else begin
        weight_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_1079_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TREADY = 1'b1;
    end else begin
        weight_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln248_fu_1079_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((ap_enable_reg_pp0_iter2 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter2 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln248_fu_1079_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accu_0_0_V_fu_1945_p2 = ($signed(add_ln700_fu_1936_p2) + $signed(sext_ln700_2_fu_1942_p1));

assign accu_0_1_V_fu_1963_p2 = ($signed(add_ln700_3_fu_1954_p2) + $signed(sext_ln700_5_fu_1960_p1));

assign accu_0_2_V_fu_1981_p2 = ($signed(add_ln700_6_fu_1972_p2) + $signed(sext_ln700_8_fu_1978_p1));

assign accu_0_3_V_fu_1999_p2 = ($signed(add_ln700_9_fu_1990_p2) + $signed(sext_ln700_11_fu_1996_p1));

assign add_ln700_10_fu_1799_p2 = ($signed(sext_ln700_10_fu_1795_p1) + $signed(sext_ln170_3_fu_1782_p1));

assign add_ln700_12_fu_2545_p2 = (zext_ln142_1_fu_2451_p1 + zext_ln142_2_fu_2460_p1);

assign add_ln700_13_fu_2555_p2 = (zext_ln700_1_fu_2551_p1 + select_ln700_fu_2438_p3);

assign add_ln700_14_fu_2561_p2 = (zext_ln142_3_fu_2469_p1 + zext_ln142_4_fu_2478_p1);

assign add_ln700_15_fu_2571_p2 = (zext_ln142_5_fu_2487_p1 + zext_ln142_6_fu_2496_p1);

assign add_ln700_16_fu_2581_p2 = (zext_ln700_3_fu_2577_p1 + zext_ln700_2_fu_2567_p1);

assign add_ln700_17_fu_2591_p2 = (zext_ln700_4_fu_2587_p1 + add_ln700_13_fu_2555_p2);

assign add_ln700_18_fu_2597_p2 = (zext_ln142_8_fu_2503_p1 + zext_ln142_9_fu_2506_p1);

assign add_ln700_19_fu_2603_p2 = (add_ln700_18_fu_2597_p2 + zext_ln142_7_fu_2500_p1);

assign add_ln700_1_fu_1676_p2 = ($signed(sext_ln700_1_fu_1672_p1) + $signed(sext_ln170_fu_1645_p1));

assign add_ln700_20_fu_2613_p2 = (zext_ln142_10_fu_2514_p1 + zext_ln142_11_fu_2523_p1);

assign add_ln700_21_fu_2623_p2 = (zext_ln142_12_fu_2532_p1 + zext_ln700_fu_2541_p1);

assign add_ln700_22_fu_2633_p2 = (zext_ln700_7_fu_2629_p1 + zext_ln700_6_fu_2619_p1);

assign add_ln700_23_fu_2639_p2 = (add_ln700_22_fu_2633_p2 + zext_ln700_5_fu_2609_p1);

assign add_ln700_24_fu_2649_p2 = (zext_ln700_8_fu_2645_p1 + add_ln700_17_fu_2591_p2);

assign add_ln700_25_fu_2767_p2 = (zext_ln142_13_fu_2673_p1 + zext_ln142_14_fu_2682_p1);

assign add_ln700_26_fu_2777_p2 = (zext_ln700_10_fu_2773_p1 + select_ln700_1_fu_2660_p3);

assign add_ln700_27_fu_2783_p2 = (zext_ln142_15_fu_2691_p1 + zext_ln142_16_fu_2700_p1);

assign add_ln700_28_fu_2793_p2 = (zext_ln142_17_fu_2709_p1 + zext_ln142_18_fu_2718_p1);

assign add_ln700_29_fu_2803_p2 = (zext_ln700_12_fu_2799_p1 + zext_ln700_11_fu_2789_p1);

assign add_ln700_30_fu_2813_p2 = (zext_ln700_13_fu_2809_p1 + add_ln700_26_fu_2777_p2);

assign add_ln700_31_fu_2819_p2 = (zext_ln142_20_fu_2725_p1 + zext_ln142_21_fu_2728_p1);

assign add_ln700_32_fu_2825_p2 = (add_ln700_31_fu_2819_p2 + zext_ln142_19_fu_2722_p1);

assign add_ln700_33_fu_2835_p2 = (zext_ln142_22_fu_2736_p1 + zext_ln142_23_fu_2745_p1);

assign add_ln700_34_fu_2845_p2 = (zext_ln142_24_fu_2754_p1 + zext_ln700_9_fu_2763_p1);

assign add_ln700_35_fu_2855_p2 = (zext_ln700_16_fu_2851_p1 + zext_ln700_15_fu_2841_p1);

assign add_ln700_36_fu_2861_p2 = (add_ln700_35_fu_2855_p2 + zext_ln700_14_fu_2831_p1);

assign add_ln700_37_fu_2871_p2 = (zext_ln700_17_fu_2867_p1 + add_ln700_30_fu_2813_p2);

assign add_ln700_38_fu_2989_p2 = (zext_ln142_25_fu_2895_p1 + zext_ln142_26_fu_2904_p1);

assign add_ln700_39_fu_2999_p2 = (zext_ln700_19_fu_2995_p1 + select_ln700_2_fu_2882_p3);

assign add_ln700_3_fu_1954_p2 = ($signed(sext_ln700_3_fu_1951_p1) + $signed(select_ln271_2_fu_1919_p3));

assign add_ln700_40_fu_3005_p2 = (zext_ln142_27_fu_2913_p1 + zext_ln142_28_fu_2922_p1);

assign add_ln700_41_fu_3015_p2 = (zext_ln142_29_fu_2931_p1 + zext_ln142_30_fu_2940_p1);

assign add_ln700_42_fu_3025_p2 = (zext_ln700_21_fu_3021_p1 + zext_ln700_20_fu_3011_p1);

assign add_ln700_43_fu_3035_p2 = (zext_ln700_22_fu_3031_p1 + add_ln700_39_fu_2999_p2);

assign add_ln700_44_fu_3041_p2 = (zext_ln142_32_fu_2947_p1 + zext_ln142_33_fu_2950_p1);

assign add_ln700_45_fu_3047_p2 = (add_ln700_44_fu_3041_p2 + zext_ln142_31_fu_2944_p1);

assign add_ln700_46_fu_3057_p2 = (zext_ln142_34_fu_2958_p1 + zext_ln142_35_fu_2967_p1);

assign add_ln700_47_fu_3067_p2 = (zext_ln142_36_fu_2976_p1 + zext_ln700_18_fu_2985_p1);

assign add_ln700_48_fu_3077_p2 = (zext_ln700_25_fu_3073_p1 + zext_ln700_24_fu_3063_p1);

assign add_ln700_49_fu_3083_p2 = (add_ln700_48_fu_3077_p2 + zext_ln700_23_fu_3053_p1);

assign add_ln700_4_fu_1717_p2 = ($signed(sext_ln700_4_fu_1713_p1) + $signed(sext_ln170_1_fu_1700_p1));

assign add_ln700_50_fu_3093_p2 = (zext_ln700_26_fu_3089_p1 + add_ln700_43_fu_3035_p2);

assign add_ln700_51_fu_3211_p2 = (zext_ln142_37_fu_3117_p1 + zext_ln142_38_fu_3126_p1);

assign add_ln700_52_fu_3221_p2 = (zext_ln700_28_fu_3217_p1 + select_ln700_3_fu_3104_p3);

assign add_ln700_53_fu_3227_p2 = (zext_ln142_39_fu_3135_p1 + zext_ln142_40_fu_3144_p1);

assign add_ln700_54_fu_3237_p2 = (zext_ln142_41_fu_3153_p1 + zext_ln142_42_fu_3162_p1);

assign add_ln700_55_fu_3247_p2 = (zext_ln700_30_fu_3243_p1 + zext_ln700_29_fu_3233_p1);

assign add_ln700_56_fu_3257_p2 = (zext_ln700_31_fu_3253_p1 + add_ln700_52_fu_3221_p2);

assign add_ln700_57_fu_3263_p2 = (zext_ln142_44_fu_3169_p1 + zext_ln142_45_fu_3172_p1);

assign add_ln700_58_fu_3269_p2 = (add_ln700_57_fu_3263_p2 + zext_ln142_43_fu_3166_p1);

assign add_ln700_59_fu_3279_p2 = (zext_ln142_46_fu_3180_p1 + zext_ln142_47_fu_3189_p1);

assign add_ln700_60_fu_3289_p2 = (zext_ln142_48_fu_3198_p1 + zext_ln700_27_fu_3207_p1);

assign add_ln700_61_fu_3299_p2 = (zext_ln700_34_fu_3295_p1 + zext_ln700_33_fu_3285_p1);

assign add_ln700_62_fu_3305_p2 = (add_ln700_61_fu_3299_p2 + zext_ln700_32_fu_3275_p1);

assign add_ln700_63_fu_3315_p2 = (zext_ln700_35_fu_3311_p1 + add_ln700_56_fu_3257_p2);

assign add_ln700_6_fu_1972_p2 = ($signed(sext_ln700_6_fu_1969_p1) + $signed(select_ln271_1_fu_1912_p3));

assign add_ln700_7_fu_1758_p2 = ($signed(sext_ln700_7_fu_1754_p1) + $signed(sext_ln170_2_fu_1741_p1));

assign add_ln700_9_fu_1990_p2 = ($signed(sext_ln700_9_fu_1987_p1) + $signed(select_ln271_fu_1905_p3));

assign add_ln700_fu_1936_p2 = ($signed(sext_ln700_fu_1933_p1) + $signed(select_ln271_3_fu_1926_p3));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state6 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op51_read_state2 == 1'b1)) | ((icmp_ln248_fu_1079_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_block_state5_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op51_read_state2 == 1'b1)) | ((icmp_ln248_fu_1079_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_block_state5_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op51_read_state2 == 1'b1)) | ((icmp_ln248_fu_1079_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op51_read_state2 == 1'b1)) | ((icmp_ln248_fu_1079_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state5_io = ((icmp_ln289_reg_3519_pp0_iter2_reg == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_485 = ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_reg_pp0_iter0_act_m_val_V_reg_1060 = 'bx;

always @ (*) begin
    ap_predicate_op51_read_state2 = ((icmp_ln252_fu_1094_p2 == 1'd1) & (icmp_ln248_fu_1079_p2 == 1'd0));
end

assign arg_V_read_assign_1_fu_1622_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1060[15:8]}};

assign arg_V_read_assign_2_fu_1649_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1060[23:16]}};

assign i_fu_1085_p2 = (i_0_reg_1049 + 17'd1);

assign icmp_ln248_fu_1079_p2 = ((i_0_reg_1049 == 17'd129600) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_1094_p2 = ((ap_sig_allocacmp_nf_assign_load_1 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln271_fu_1468_p2 = ((sf_1_fu_258 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln289_fu_1594_p2 = ((sf_fu_1588_p2 == 32'd9) ? 1'b1 : 1'b0);

assign icmp_ln301_fu_1874_p2 = ((nf_fu_1868_p2 == 32'd16) ? 1'b1 : 1'b0);

assign icmp_ln321_1_fu_1168_p2 = ((trunc_ln321_fu_1158_p1 == 4'd6) ? 1'b1 : 1'b0);

assign icmp_ln321_2_fu_1174_p2 = ((trunc_ln321_fu_1158_p1 == 4'd5) ? 1'b1 : 1'b0);

assign icmp_ln321_3_fu_1180_p2 = ((trunc_ln321_fu_1158_p1 == 4'd4) ? 1'b1 : 1'b0);

assign icmp_ln321_4_fu_1186_p2 = ((trunc_ln321_fu_1158_p1 == 4'd3) ? 1'b1 : 1'b0);

assign icmp_ln321_5_fu_1192_p2 = ((trunc_ln321_fu_1158_p1 == 4'd2) ? 1'b1 : 1'b0);

assign icmp_ln321_6_fu_1198_p2 = ((trunc_ln321_fu_1158_p1 == 4'd1) ? 1'b1 : 1'b0);

assign icmp_ln321_7_fu_1204_p2 = ((trunc_ln321_fu_1158_p1 == 4'd0) ? 1'b1 : 1'b0);

assign icmp_ln321_fu_1162_p2 = ((trunc_ln321_fu_1158_p1 == 4'd7) ? 1'b1 : 1'b0);

assign icmp_ln899_10_fu_2103_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_53_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_11_fu_2109_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_52_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_12_fu_2115_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_51_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_13_fu_2121_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_50_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_14_fu_2127_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_41_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_15_fu_2133_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_40_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_16_fu_2139_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_35_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_17_fu_2145_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_34_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_18_fu_2151_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_33_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_19_fu_2157_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_32_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_1_fu_2031_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_54_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_20_fu_2163_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_31_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_21_fu_2169_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_30_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_22_fu_2181_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_29_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_23_fu_2193_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_28_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_24_fu_2205_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_39_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_25_fu_2211_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_38_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_26_fu_2217_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_37_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_27_fu_2223_p2 = (($signed(accu_0_1_V_fu_1963_p2) < $signed(threshs_m_thresholds_36_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_28_fu_2229_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_27_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_29_fu_2235_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_26_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_2_fu_2037_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_49_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_30_fu_2241_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_21_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_31_fu_2247_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_20_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_32_fu_2253_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_19_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_33_fu_2259_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_18_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_34_fu_2265_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_17_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_35_fu_2271_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_16_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_36_fu_2283_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_15_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_37_fu_2295_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_14_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_38_fu_2307_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_25_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_39_fu_2313_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_24_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_3_fu_2043_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_48_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_40_fu_2319_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_23_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_41_fu_2325_p2 = (($signed(accu_0_2_V_fu_1981_p2) < $signed(threshs_m_thresholds_22_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_42_fu_2331_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_13_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_43_fu_2337_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_12_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_44_fu_2343_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_7_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_45_fu_2349_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_6_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_46_fu_2355_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_5_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_47_fu_2361_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_4_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_48_fu_2367_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_3_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_49_fu_2373_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_2_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_4_fu_2049_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_47_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_50_fu_2385_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_1_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_51_fu_2397_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_52_fu_2409_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_11_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_53_fu_2415_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_10_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_54_fu_2421_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_9_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_55_fu_2427_p2 = (($signed(accu_0_3_V_fu_1999_p2) < $signed(threshs_m_thresholds_8_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_5_fu_2055_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_46_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_6_fu_2061_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_45_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_7_fu_2067_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_44_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_8_fu_2079_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_43_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_9_fu_2091_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_42_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_fu_2025_p2 = (($signed(accu_0_0_V_fu_1945_p2) < $signed(threshs_m_thresholds_55_q0)) ? 1'b1 : 1'b0);

assign inElem_V_fu_1134_p10 = sf_1_fu_258[3:0];

assign inputBuf_8_V_11_fu_1284_p3 = ((or_ln321_6_fu_1246_p2[0:0] === 1'b1) ? select_ln321_2_fu_1276_p3 : inputBuf_8_V_8_fu_294);

assign inputBuf_8_V_12_fu_1308_p3 = ((or_ln321_4_fu_1234_p2[0:0] === 1'b1) ? inputBuf_8_V_3_fu_290 : select_ln321_5_fu_1300_p3);

assign inputBuf_8_V_13_fu_1332_p3 = ((or_ln321_4_fu_1234_p2[0:0] === 1'b1) ? inputBuf_8_V_5_fu_286 : select_ln321_8_fu_1324_p3);

assign inputBuf_8_V_14_fu_1348_p3 = ((or_ln321_4_fu_1234_p2[0:0] === 1'b1) ? inputBuf_8_V_7_fu_282 : select_ln321_10_fu_1340_p3);

assign inputBuf_8_V_15_fu_1372_p3 = ((or_ln321_4_fu_1234_p2[0:0] === 1'b1) ? select_ln321_13_fu_1364_p3 : inputBuf_8_V_6_fu_278);

assign inputBuf_8_V_16_fu_1388_p3 = ((or_ln321_fu_1210_p2[0:0] === 1'b1) ? inputBuf_8_V_4_fu_274 : select_ln321_15_fu_1380_p3);

assign inputBuf_8_V_17_fu_1396_p3 = ((icmp_ln321_6_fu_1198_p2[0:0] === 1'b1) ? in_V_V_TDATA : inputBuf_8_V_2_fu_270);

assign inputBuf_8_V_18_fu_1404_p3 = ((icmp_ln321_7_fu_1204_p2[0:0] === 1'b1) ? inputBuf_8_V_2_fu_270 : inputBuf_8_V_17_fu_1396_p3);

assign inputBuf_8_V_19_fu_1412_p3 = ((icmp_ln321_7_fu_1204_p2[0:0] === 1'b1) ? in_V_V_TDATA : inputBuf_8_V_1_fu_266);

assign inputBuf_8_V_fu_1252_p3 = ((or_ln321_6_fu_1246_p2[0:0] === 1'b1) ? inputBuf_8_V_9_fu_298 : in_V_V_TDATA);

assign mul_ln1352_10_fu_1776_p0 = sext_ln215_3_fu_1635_p1;

assign mul_ln1352_11_fu_1789_p0 = sext_ln215_5_fu_1662_p1;

assign mul_ln1352_1_fu_1639_p0 = sext_ln215_3_fu_1635_p1;

assign mul_ln1352_2_fu_1666_p0 = sext_ln215_5_fu_1662_p1;

assign mul_ln1352_3_fu_1685_p0 = sext_ln215_1_fu_1612_p1;

assign mul_ln1352_4_fu_1694_p0 = sext_ln215_3_fu_1635_p1;

assign mul_ln1352_5_fu_1707_p0 = sext_ln215_5_fu_1662_p1;

assign mul_ln1352_6_fu_1726_p0 = sext_ln215_1_fu_1612_p1;

assign mul_ln1352_7_fu_1735_p0 = sext_ln215_3_fu_1635_p1;

assign mul_ln1352_8_fu_1748_p0 = sext_ln215_5_fu_1662_p1;

assign mul_ln1352_9_fu_1767_p0 = sext_ln215_1_fu_1612_p1;

assign mul_ln1352_fu_1616_p0 = sext_ln215_1_fu_1612_p1;

assign nf_fu_1868_p2 = (nf_assign_fu_262 + 32'd1);

assign or_ln321_1_fu_1216_p2 = (icmp_ln321_5_fu_1192_p2 | icmp_ln321_4_fu_1186_p2);

assign or_ln321_2_fu_1222_p2 = (icmp_ln321_3_fu_1180_p2 | icmp_ln321_2_fu_1174_p2);

assign or_ln321_3_fu_1228_p2 = (icmp_ln321_fu_1162_p2 | icmp_ln321_1_fu_1168_p2);

assign or_ln321_4_fu_1234_p2 = (or_ln321_fu_1210_p2 | or_ln321_1_fu_1216_p2);

assign or_ln321_5_fu_1240_p2 = (or_ln321_3_fu_1228_p2 | or_ln321_2_fu_1222_p2);

assign or_ln321_6_fu_1246_p2 = (or_ln321_5_fu_1240_p2 | or_ln321_4_fu_1234_p2);

assign or_ln321_fu_1210_p2 = (icmp_ln321_7_fu_1204_p2 | icmp_ln321_6_fu_1198_p2);

assign out_V_V_TDATA = {{{{add_ln700_63_fu_3315_p2}, {add_ln700_50_fu_3093_p2}}, {add_ln700_37_fu_2871_p2}}, {add_ln700_24_fu_2649_p2}};

assign select_ln271_1_fu_1912_p3 = ((icmp_ln271_reg_3451_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_2_0_fu_250);

assign select_ln271_2_fu_1919_p3 = ((icmp_ln271_reg_3451_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_1_0_fu_246);

assign select_ln271_3_fu_1926_p3 = ((icmp_ln271_reg_3451_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_0_0_fu_242);

assign select_ln271_fu_1905_p3 = ((icmp_ln271_reg_3451_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_3_0_fu_254);

assign select_ln301_fu_1880_p3 = ((icmp_ln301_fu_1874_p2[0:0] === 1'b1) ? 32'd0 : nf_fu_1868_p2);

assign select_ln321_10_fu_1340_p3 = ((icmp_ln321_3_fu_1180_p2[0:0] === 1'b1) ? in_V_V_TDATA : inputBuf_8_V_7_fu_282);

assign select_ln321_12_fu_1356_p3 = ((icmp_ln321_5_fu_1192_p2[0:0] === 1'b1) ? inputBuf_8_V_6_fu_278 : in_V_V_TDATA);

assign select_ln321_13_fu_1364_p3 = ((or_ln321_fu_1210_p2[0:0] === 1'b1) ? inputBuf_8_V_6_fu_278 : select_ln321_12_fu_1356_p3);

assign select_ln321_15_fu_1380_p3 = ((icmp_ln321_5_fu_1192_p2[0:0] === 1'b1) ? in_V_V_TDATA : inputBuf_8_V_4_fu_274);

assign select_ln321_1_fu_1268_p3 = ((or_ln321_2_fu_1222_p2[0:0] === 1'b1) ? inputBuf_8_V_8_fu_294 : select_ln321_fu_1260_p3);

assign select_ln321_2_fu_1276_p3 = ((or_ln321_4_fu_1234_p2[0:0] === 1'b1) ? inputBuf_8_V_8_fu_294 : select_ln321_1_fu_1268_p3);

assign select_ln321_4_fu_1292_p3 = ((icmp_ln321_1_fu_1168_p2[0:0] === 1'b1) ? in_V_V_TDATA : inputBuf_8_V_3_fu_290);

assign select_ln321_5_fu_1300_p3 = ((or_ln321_2_fu_1222_p2[0:0] === 1'b1) ? inputBuf_8_V_3_fu_290 : select_ln321_4_fu_1292_p3);

assign select_ln321_7_fu_1316_p3 = ((icmp_ln321_3_fu_1180_p2[0:0] === 1'b1) ? inputBuf_8_V_5_fu_286 : in_V_V_TDATA);

assign select_ln321_8_fu_1324_p3 = ((or_ln321_2_fu_1222_p2[0:0] === 1'b1) ? select_ln321_7_fu_1316_p3 : inputBuf_8_V_5_fu_286);

assign select_ln321_fu_1260_p3 = ((icmp_ln321_1_fu_1168_p2[0:0] === 1'b1) ? inputBuf_8_V_8_fu_294 : in_V_V_TDATA);

assign select_ln700_1_fu_2660_p3 = ((xor_ln899_14_fu_2655_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign select_ln700_2_fu_2882_p3 = ((xor_ln899_28_fu_2877_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign select_ln700_3_fu_3104_p3 = ((xor_ln899_42_fu_3099_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign select_ln700_fu_2438_p3 = ((xor_ln899_fu_2433_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign sext_ln170_1_fu_1700_p1 = mul_ln1352_4_fu_1694_p2;

assign sext_ln170_2_fu_1741_p1 = mul_ln1352_7_fu_1735_p2;

assign sext_ln170_3_fu_1782_p1 = mul_ln1352_10_fu_1776_p2;

assign sext_ln170_fu_1645_p1 = mul_ln1352_1_fu_1639_p2;

assign sext_ln215_1_fu_1612_p1 = $signed(trunc_ln647_1_fu_1605_p1);

assign sext_ln215_3_fu_1635_p1 = $signed(arg_V_read_assign_1_fu_1622_p4);

assign sext_ln215_5_fu_1662_p1 = $signed(arg_V_read_assign_2_fu_1649_p4);

assign sext_ln700_10_fu_1795_p1 = mul_ln1352_11_fu_1789_p2;

assign sext_ln700_11_fu_1996_p1 = $signed(add_ln700_10_reg_3558);

assign sext_ln700_1_fu_1672_p1 = mul_ln1352_2_fu_1666_p2;

assign sext_ln700_2_fu_1942_p1 = $signed(add_ln700_1_reg_3528);

assign sext_ln700_3_fu_1951_p1 = mul_ln1352_3_reg_3533;

assign sext_ln700_4_fu_1713_p1 = mul_ln1352_5_fu_1707_p2;

assign sext_ln700_5_fu_1960_p1 = $signed(add_ln700_4_reg_3538);

assign sext_ln700_6_fu_1969_p1 = mul_ln1352_6_reg_3543;

assign sext_ln700_7_fu_1754_p1 = mul_ln1352_8_fu_1748_p2;

assign sext_ln700_8_fu_1978_p1 = $signed(add_ln700_7_reg_3548);

assign sext_ln700_9_fu_1987_p1 = mul_ln1352_9_reg_3553;

assign sext_ln700_fu_1933_p1 = mul_ln1352_reg_3523;

assign sf_fu_1588_p2 = (32'd1 + sf_1_fu_258);

assign threshs_m_thresholds_10_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_11_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_12_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_13_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_14_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_15_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_16_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_17_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_18_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_19_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_1_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_20_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_21_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_22_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_23_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_24_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_25_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_26_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_27_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_28_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_29_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_2_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_30_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_31_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_32_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_33_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_34_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_35_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_36_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_37_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_38_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_39_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_3_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_40_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_41_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_42_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_43_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_44_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_45_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_46_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_47_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_48_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_49_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_4_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_50_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_51_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_52_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_53_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_54_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_55_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_5_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_6_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_7_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_8_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_9_address0 = zext_ln142_fu_1808_p1;

assign threshs_m_thresholds_address0 = zext_ln142_fu_1808_p1;

assign trunc_ln321_fu_1158_p1 = sf_1_fu_258[3:0];

assign trunc_ln647_1_fu_1605_p1 = ap_phi_reg_pp0_iter1_act_m_val_V_reg_1060[7:0];

assign trunc_ln647_fu_1474_p1 = weight_V_V_TDATA[3:0];

assign xor_ln899_10_fu_2509_p2 = (icmp_ln899_10_reg_3893 ^ 1'd1);

assign xor_ln899_11_fu_2518_p2 = (icmp_ln899_11_reg_3898 ^ 1'd1);

assign xor_ln899_12_fu_2527_p2 = (icmp_ln899_12_reg_3903 ^ 1'd1);

assign xor_ln899_13_fu_2536_p2 = (icmp_ln899_13_reg_3908 ^ 1'd1);

assign xor_ln899_14_fu_2655_p2 = (icmp_ln899_14_reg_3913 ^ 1'd1);

assign xor_ln899_15_fu_2668_p2 = (icmp_ln899_15_reg_3918 ^ 1'd1);

assign xor_ln899_16_fu_2677_p2 = (icmp_ln899_16_reg_3923 ^ 1'd1);

assign xor_ln899_17_fu_2686_p2 = (icmp_ln899_17_reg_3928 ^ 1'd1);

assign xor_ln899_18_fu_2695_p2 = (icmp_ln899_18_reg_3933 ^ 1'd1);

assign xor_ln899_19_fu_2704_p2 = (icmp_ln899_19_reg_3938 ^ 1'd1);

assign xor_ln899_1_fu_2446_p2 = (icmp_ln899_1_reg_3848 ^ 1'd1);

assign xor_ln899_20_fu_2713_p2 = (icmp_ln899_20_reg_3943 ^ 1'd1);

assign xor_ln899_21_fu_2175_p2 = (icmp_ln899_21_fu_2169_p2 ^ 1'd1);

assign xor_ln899_22_fu_2187_p2 = (icmp_ln899_22_fu_2181_p2 ^ 1'd1);

assign xor_ln899_23_fu_2199_p2 = (icmp_ln899_23_fu_2193_p2 ^ 1'd1);

assign xor_ln899_24_fu_2731_p2 = (icmp_ln899_24_reg_3963 ^ 1'd1);

assign xor_ln899_25_fu_2740_p2 = (icmp_ln899_25_reg_3968 ^ 1'd1);

assign xor_ln899_26_fu_2749_p2 = (icmp_ln899_26_reg_3973 ^ 1'd1);

assign xor_ln899_27_fu_2758_p2 = (icmp_ln899_27_reg_3978 ^ 1'd1);

assign xor_ln899_28_fu_2877_p2 = (icmp_ln899_28_reg_3983 ^ 1'd1);

assign xor_ln899_29_fu_2890_p2 = (icmp_ln899_29_reg_3988 ^ 1'd1);

assign xor_ln899_2_fu_2455_p2 = (icmp_ln899_2_reg_3853 ^ 1'd1);

assign xor_ln899_30_fu_2899_p2 = (icmp_ln899_30_reg_3993 ^ 1'd1);

assign xor_ln899_31_fu_2908_p2 = (icmp_ln899_31_reg_3998 ^ 1'd1);

assign xor_ln899_32_fu_2917_p2 = (icmp_ln899_32_reg_4003 ^ 1'd1);

assign xor_ln899_33_fu_2926_p2 = (icmp_ln899_33_reg_4008 ^ 1'd1);

assign xor_ln899_34_fu_2935_p2 = (icmp_ln899_34_reg_4013 ^ 1'd1);

assign xor_ln899_35_fu_2277_p2 = (icmp_ln899_35_fu_2271_p2 ^ 1'd1);

assign xor_ln899_36_fu_2289_p2 = (icmp_ln899_36_fu_2283_p2 ^ 1'd1);

assign xor_ln899_37_fu_2301_p2 = (icmp_ln899_37_fu_2295_p2 ^ 1'd1);

assign xor_ln899_38_fu_2953_p2 = (icmp_ln899_38_reg_4033 ^ 1'd1);

assign xor_ln899_39_fu_2962_p2 = (icmp_ln899_39_reg_4038 ^ 1'd1);

assign xor_ln899_3_fu_2464_p2 = (icmp_ln899_3_reg_3858 ^ 1'd1);

assign xor_ln899_40_fu_2971_p2 = (icmp_ln899_40_reg_4043 ^ 1'd1);

assign xor_ln899_41_fu_2980_p2 = (icmp_ln899_41_reg_4048 ^ 1'd1);

assign xor_ln899_42_fu_3099_p2 = (icmp_ln899_42_reg_4053 ^ 1'd1);

assign xor_ln899_43_fu_3112_p2 = (icmp_ln899_43_reg_4058 ^ 1'd1);

assign xor_ln899_44_fu_3121_p2 = (icmp_ln899_44_reg_4063 ^ 1'd1);

assign xor_ln899_45_fu_3130_p2 = (icmp_ln899_45_reg_4068 ^ 1'd1);

assign xor_ln899_46_fu_3139_p2 = (icmp_ln899_46_reg_4073 ^ 1'd1);

assign xor_ln899_47_fu_3148_p2 = (icmp_ln899_47_reg_4078 ^ 1'd1);

assign xor_ln899_48_fu_3157_p2 = (icmp_ln899_48_reg_4083 ^ 1'd1);

assign xor_ln899_49_fu_2379_p2 = (icmp_ln899_49_fu_2373_p2 ^ 1'd1);

assign xor_ln899_4_fu_2473_p2 = (icmp_ln899_4_reg_3863 ^ 1'd1);

assign xor_ln899_50_fu_2391_p2 = (icmp_ln899_50_fu_2385_p2 ^ 1'd1);

assign xor_ln899_51_fu_2403_p2 = (icmp_ln899_51_fu_2397_p2 ^ 1'd1);

assign xor_ln899_52_fu_3175_p2 = (icmp_ln899_52_reg_4103 ^ 1'd1);

assign xor_ln899_53_fu_3184_p2 = (icmp_ln899_53_reg_4108 ^ 1'd1);

assign xor_ln899_54_fu_3193_p2 = (icmp_ln899_54_reg_4113 ^ 1'd1);

assign xor_ln899_55_fu_3202_p2 = (icmp_ln899_55_reg_4118 ^ 1'd1);

assign xor_ln899_5_fu_2482_p2 = (icmp_ln899_5_reg_3868 ^ 1'd1);

assign xor_ln899_6_fu_2491_p2 = (icmp_ln899_6_reg_3873 ^ 1'd1);

assign xor_ln899_7_fu_2073_p2 = (icmp_ln899_7_fu_2067_p2 ^ 1'd1);

assign xor_ln899_8_fu_2085_p2 = (icmp_ln899_8_fu_2079_p2 ^ 1'd1);

assign xor_ln899_9_fu_2097_p2 = (icmp_ln899_9_fu_2091_p2 ^ 1'd1);

assign xor_ln899_fu_2433_p2 = (icmp_ln899_reg_3843 ^ 1'd1);

assign zext_ln142_10_fu_2514_p1 = xor_ln899_10_fu_2509_p2;

assign zext_ln142_11_fu_2523_p1 = xor_ln899_11_fu_2518_p2;

assign zext_ln142_12_fu_2532_p1 = xor_ln899_12_fu_2527_p2;

assign zext_ln142_13_fu_2673_p1 = xor_ln899_15_fu_2668_p2;

assign zext_ln142_14_fu_2682_p1 = xor_ln899_16_fu_2677_p2;

assign zext_ln142_15_fu_2691_p1 = xor_ln899_17_fu_2686_p2;

assign zext_ln142_16_fu_2700_p1 = xor_ln899_18_fu_2695_p2;

assign zext_ln142_17_fu_2709_p1 = xor_ln899_19_fu_2704_p2;

assign zext_ln142_18_fu_2718_p1 = xor_ln899_20_fu_2713_p2;

assign zext_ln142_19_fu_2722_p1 = xor_ln899_21_reg_3948;

assign zext_ln142_1_fu_2451_p1 = xor_ln899_1_fu_2446_p2;

assign zext_ln142_20_fu_2725_p1 = xor_ln899_22_reg_3953;

assign zext_ln142_21_fu_2728_p1 = xor_ln899_23_reg_3958;

assign zext_ln142_22_fu_2736_p1 = xor_ln899_24_fu_2731_p2;

assign zext_ln142_23_fu_2745_p1 = xor_ln899_25_fu_2740_p2;

assign zext_ln142_24_fu_2754_p1 = xor_ln899_26_fu_2749_p2;

assign zext_ln142_25_fu_2895_p1 = xor_ln899_29_fu_2890_p2;

assign zext_ln142_26_fu_2904_p1 = xor_ln899_30_fu_2899_p2;

assign zext_ln142_27_fu_2913_p1 = xor_ln899_31_fu_2908_p2;

assign zext_ln142_28_fu_2922_p1 = xor_ln899_32_fu_2917_p2;

assign zext_ln142_29_fu_2931_p1 = xor_ln899_33_fu_2926_p2;

assign zext_ln142_2_fu_2460_p1 = xor_ln899_2_fu_2455_p2;

assign zext_ln142_30_fu_2940_p1 = xor_ln899_34_fu_2935_p2;

assign zext_ln142_31_fu_2944_p1 = xor_ln899_35_reg_4018;

assign zext_ln142_32_fu_2947_p1 = xor_ln899_36_reg_4023;

assign zext_ln142_33_fu_2950_p1 = xor_ln899_37_reg_4028;

assign zext_ln142_34_fu_2958_p1 = xor_ln899_38_fu_2953_p2;

assign zext_ln142_35_fu_2967_p1 = xor_ln899_39_fu_2962_p2;

assign zext_ln142_36_fu_2976_p1 = xor_ln899_40_fu_2971_p2;

assign zext_ln142_37_fu_3117_p1 = xor_ln899_43_fu_3112_p2;

assign zext_ln142_38_fu_3126_p1 = xor_ln899_44_fu_3121_p2;

assign zext_ln142_39_fu_3135_p1 = xor_ln899_45_fu_3130_p2;

assign zext_ln142_3_fu_2469_p1 = xor_ln899_3_fu_2464_p2;

assign zext_ln142_40_fu_3144_p1 = xor_ln899_46_fu_3139_p2;

assign zext_ln142_41_fu_3153_p1 = xor_ln899_47_fu_3148_p2;

assign zext_ln142_42_fu_3162_p1 = xor_ln899_48_fu_3157_p2;

assign zext_ln142_43_fu_3166_p1 = xor_ln899_49_reg_4088;

assign zext_ln142_44_fu_3169_p1 = xor_ln899_50_reg_4093;

assign zext_ln142_45_fu_3172_p1 = xor_ln899_51_reg_4098;

assign zext_ln142_46_fu_3180_p1 = xor_ln899_52_fu_3175_p2;

assign zext_ln142_47_fu_3189_p1 = xor_ln899_53_fu_3184_p2;

assign zext_ln142_48_fu_3198_p1 = xor_ln899_54_fu_3193_p2;

assign zext_ln142_4_fu_2478_p1 = xor_ln899_4_fu_2473_p2;

assign zext_ln142_5_fu_2487_p1 = xor_ln899_5_fu_2482_p2;

assign zext_ln142_6_fu_2496_p1 = xor_ln899_6_fu_2491_p2;

assign zext_ln142_7_fu_2500_p1 = xor_ln899_7_reg_3878;

assign zext_ln142_8_fu_2503_p1 = xor_ln899_8_reg_3883;

assign zext_ln142_9_fu_2506_p1 = xor_ln899_9_reg_3888;

assign zext_ln142_fu_1808_p1 = nf_assign_fu_262;

assign zext_ln700_10_fu_2773_p1 = add_ln700_25_fu_2767_p2;

assign zext_ln700_11_fu_2789_p1 = add_ln700_27_fu_2783_p2;

assign zext_ln700_12_fu_2799_p1 = add_ln700_28_fu_2793_p2;

assign zext_ln700_13_fu_2809_p1 = add_ln700_29_fu_2803_p2;

assign zext_ln700_14_fu_2831_p1 = add_ln700_32_fu_2825_p2;

assign zext_ln700_15_fu_2841_p1 = add_ln700_33_fu_2835_p2;

assign zext_ln700_16_fu_2851_p1 = add_ln700_34_fu_2845_p2;

assign zext_ln700_17_fu_2867_p1 = add_ln700_36_fu_2861_p2;

assign zext_ln700_18_fu_2985_p1 = xor_ln899_41_fu_2980_p2;

assign zext_ln700_19_fu_2995_p1 = add_ln700_38_fu_2989_p2;

assign zext_ln700_1_fu_2551_p1 = add_ln700_12_fu_2545_p2;

assign zext_ln700_20_fu_3011_p1 = add_ln700_40_fu_3005_p2;

assign zext_ln700_21_fu_3021_p1 = add_ln700_41_fu_3015_p2;

assign zext_ln700_22_fu_3031_p1 = add_ln700_42_fu_3025_p2;

assign zext_ln700_23_fu_3053_p1 = add_ln700_45_fu_3047_p2;

assign zext_ln700_24_fu_3063_p1 = add_ln700_46_fu_3057_p2;

assign zext_ln700_25_fu_3073_p1 = add_ln700_47_fu_3067_p2;

assign zext_ln700_26_fu_3089_p1 = add_ln700_49_fu_3083_p2;

assign zext_ln700_27_fu_3207_p1 = xor_ln899_55_fu_3202_p2;

assign zext_ln700_28_fu_3217_p1 = add_ln700_51_fu_3211_p2;

assign zext_ln700_29_fu_3233_p1 = add_ln700_53_fu_3227_p2;

assign zext_ln700_2_fu_2567_p1 = add_ln700_14_fu_2561_p2;

assign zext_ln700_30_fu_3243_p1 = add_ln700_54_fu_3237_p2;

assign zext_ln700_31_fu_3253_p1 = add_ln700_55_fu_3247_p2;

assign zext_ln700_32_fu_3275_p1 = add_ln700_58_fu_3269_p2;

assign zext_ln700_33_fu_3285_p1 = add_ln700_59_fu_3279_p2;

assign zext_ln700_34_fu_3295_p1 = add_ln700_60_fu_3289_p2;

assign zext_ln700_35_fu_3311_p1 = add_ln700_62_fu_3305_p2;

assign zext_ln700_3_fu_2577_p1 = add_ln700_15_fu_2571_p2;

assign zext_ln700_4_fu_2587_p1 = add_ln700_16_fu_2581_p2;

assign zext_ln700_5_fu_2609_p1 = add_ln700_19_fu_2603_p2;

assign zext_ln700_6_fu_2619_p1 = add_ln700_20_fu_2613_p2;

assign zext_ln700_7_fu_2629_p1 = add_ln700_21_fu_2623_p2;

assign zext_ln700_8_fu_2645_p1 = add_ln700_23_fu_2639_p2;

assign zext_ln700_9_fu_2763_p1 = xor_ln899_27_fu_2758_p2;

assign zext_ln700_fu_2541_p1 = xor_ln899_13_fu_2536_p2;

endmodule //StreamingFCLayer_Batch_2_Matrix_Vector_Activa
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Acttde.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Acttde_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Acttde_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Acttde(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Acttde_rom StreamingFCLayer_Batch_4_Matrix_Vector_Acttde_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcg8j.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_Batcg8j_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcg8j_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_Batcg8j(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_Batcg8j_rom Thresholding_Batch_1_Thresholding_Batcg8j_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActBew.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActBew_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActBew_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActBew(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActBew_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActBew_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbCo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcbCo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbCo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcbCo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcbCo_rom Thresholding_Batch_0_Thresholding_BatcbCo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_BatcfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_BatcfYi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_BatcfYi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_BatcfYi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_BatcfYi_rom Thresholding_Batch_2_Thresholding_BatcfYi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/be37/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActOgC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActOgC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActOgC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActOgC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActOgC_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActOgC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcHfu.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcHfu_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcHfu_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcHfu(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcHfu_rom Thresholding_Batch_0_Thresholding_BatcHfu_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ce70/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcibs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcibs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 4;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcibs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcibs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd4;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcibs_rom Thresholding_Batch_0_Thresholding_Batcibs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actcud.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actcud_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actcud_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actcud(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actcud_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actcud_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/cd9c/hdl/verilog/StreamingFCLayer_Batch_0_Matrix_Vector_Activa.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingFCLayer_Batch_0_Matrix_Vector_Activa (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY,
        weight_V_V_TDATA,
        weight_V_V_TVALID,
        weight_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [7:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [95:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;
input  [31:0] weight_V_V_TDATA;
input   weight_V_V_TVALID;
output   weight_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;
reg weight_V_V_TREADY;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln248_fu_4769_p2;
wire   [0:0] icmp_ln252_fu_4784_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln289_reg_15104;
reg    weight_V_V_TDATA_blk_n;
reg   [20:0] i_0_reg_3589;
reg    ap_predicate_op1183_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [20:0] i_fu_4775_p2;
wire   [7:0] inElem_V_1_fu_6525_p578;
wire   [9:0] trunc_ln321_fu_7683_p1;
wire   [0:0] icmp_ln271_fu_10570_p2;
reg   [0:0] icmp_ln271_reg_15056;
wire   [3:0] trunc_ln647_fu_10576_p1;
reg  signed [3:0] trunc_ln647_reg_15064;
reg  signed [3:0] p_Result_1_0_1_reg_15069;
reg  signed [3:0] p_Result_1_1_reg_15074;
reg  signed [3:0] p_Result_1_1_1_reg_15079;
reg  signed [3:0] p_Result_1_2_reg_15084;
reg  signed [3:0] p_Result_1_2_1_reg_15089;
reg  signed [3:0] p_Result_1_3_reg_15094;
reg  signed [3:0] p_Result_1_3_1_reg_15099;
wire   [0:0] icmp_ln289_fu_10656_p2;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
wire   [7:0] ap_phi_reg_pp0_iter0_act_m_val_V_reg_3600;
reg   [7:0] ap_phi_reg_pp0_iter1_act_m_val_V_reg_3600;
reg   [23:0] accu_0_0_V_1_fu_1242;
wire   [23:0] accu_0_0_V_fu_10765_p2;
reg   [23:0] accu_0_1_V_1_fu_1246;
wire   [23:0] accu_0_1_V_fu_10807_p2;
reg   [23:0] accu_0_2_V_1_fu_1250;
wire   [23:0] accu_0_2_V_fu_10849_p2;
reg   [23:0] accu_0_3_V_1_fu_1254;
wire   [23:0] accu_0_3_V_fu_10891_p2;
reg   [31:0] sf_1_fu_1258;
wire   [31:0] sf_fu_10650_p2;
reg   [7:0] tmp_V_fu_1262;
reg   [7:0] tmp_V_1_fu_1266;
reg   [7:0] tmp_V_2_fu_1270;
reg   [7:0] tmp_V_4_fu_1274;
reg   [7:0] tmp_V_5_fu_1278;
reg   [7:0] tmp_V_6_fu_1282;
reg   [7:0] tmp_V_7_fu_1286;
reg   [7:0] tmp_V_8_fu_1290;
reg   [7:0] tmp_V_9_fu_1294;
reg   [7:0] tmp_V_10_fu_1298;
reg   [7:0] tmp_V_11_fu_1302;
reg   [7:0] tmp_V_12_fu_1306;
reg   [7:0] tmp_V_13_fu_1310;
reg   [7:0] tmp_V_14_fu_1314;
reg   [7:0] tmp_V_15_fu_1318;
reg   [7:0] tmp_V_16_fu_1322;
reg   [7:0] tmp_V_17_fu_1326;
reg   [7:0] tmp_V_18_fu_1330;
reg   [7:0] tmp_V_19_fu_1334;
reg   [7:0] tmp_V_20_fu_1338;
reg   [7:0] tmp_V_21_fu_1342;
reg   [7:0] tmp_V_22_fu_1346;
reg   [7:0] tmp_V_23_fu_1350;
reg   [7:0] tmp_V_24_fu_1354;
reg   [7:0] tmp_V_25_fu_1358;
reg   [7:0] tmp_V_26_fu_1362;
reg   [7:0] tmp_V_27_fu_1366;
reg   [7:0] tmp_V_28_fu_1370;
reg   [7:0] tmp_V_29_fu_1374;
reg   [7:0] tmp_V_30_fu_1378;
reg   [7:0] tmp_V_31_fu_1382;
reg   [7:0] tmp_V_32_fu_1386;
reg   [7:0] tmp_V_33_fu_1390;
reg   [7:0] tmp_V_34_fu_1394;
reg   [7:0] tmp_V_35_fu_1398;
reg   [7:0] tmp_V_36_fu_1402;
reg   [7:0] tmp_V_37_fu_1406;
reg   [7:0] tmp_V_38_fu_1410;
reg   [7:0] tmp_V_39_fu_1414;
reg   [7:0] tmp_V_40_fu_1418;
reg   [7:0] tmp_V_41_fu_1422;
reg   [7:0] tmp_V_42_fu_1426;
reg   [7:0] tmp_V_43_fu_1430;
reg   [7:0] tmp_V_44_fu_1434;
reg   [7:0] tmp_V_45_fu_1438;
reg   [7:0] tmp_V_46_fu_1442;
reg   [7:0] tmp_V_47_fu_1446;
reg   [7:0] tmp_V_48_fu_1450;
reg   [7:0] tmp_V_49_fu_1454;
reg   [7:0] tmp_V_50_fu_1458;
reg   [7:0] tmp_V_51_fu_1462;
reg   [7:0] tmp_V_52_fu_1466;
reg   [7:0] tmp_V_53_fu_1470;
reg   [7:0] tmp_V_54_fu_1474;
reg   [7:0] tmp_V_55_fu_1478;
reg   [7:0] tmp_V_56_fu_1482;
reg   [7:0] tmp_V_57_fu_1486;
reg   [7:0] tmp_V_58_fu_1490;
reg   [7:0] tmp_V_59_fu_1494;
reg   [7:0] tmp_V_60_fu_1498;
reg   [7:0] tmp_V_61_fu_1502;
reg   [7:0] tmp_V_62_fu_1506;
reg   [7:0] tmp_V_63_fu_1510;
reg   [7:0] tmp_V_64_fu_1514;
reg   [7:0] tmp_V_65_fu_1518;
reg   [7:0] tmp_V_66_fu_1522;
reg   [7:0] tmp_V_67_fu_1526;
reg   [7:0] tmp_V_68_fu_1530;
reg   [7:0] tmp_V_69_fu_1534;
reg   [7:0] tmp_V_70_fu_1538;
reg   [7:0] tmp_V_71_fu_1542;
reg   [7:0] tmp_V_72_fu_1546;
reg   [7:0] tmp_V_73_fu_1550;
reg   [7:0] tmp_V_74_fu_1554;
reg   [7:0] tmp_V_75_fu_1558;
reg   [7:0] tmp_V_76_fu_1562;
reg   [7:0] tmp_V_77_fu_1566;
reg   [7:0] tmp_V_78_fu_1570;
reg   [7:0] tmp_V_79_fu_1574;
reg   [7:0] tmp_V_80_fu_1578;
reg   [7:0] tmp_V_81_fu_1582;
reg   [7:0] tmp_V_82_fu_1586;
reg   [7:0] tmp_V_83_fu_1590;
reg   [7:0] tmp_V_84_fu_1594;
reg   [7:0] tmp_V_85_fu_1598;
reg   [7:0] tmp_V_86_fu_1602;
reg   [7:0] tmp_V_87_fu_1606;
reg   [7:0] tmp_V_88_fu_1610;
reg   [7:0] tmp_V_89_fu_1614;
reg   [7:0] tmp_V_90_fu_1618;
reg   [7:0] tmp_V_91_fu_1622;
reg   [7:0] tmp_V_92_fu_1626;
reg   [7:0] tmp_V_93_fu_1630;
reg   [7:0] tmp_V_94_fu_1634;
reg   [7:0] tmp_V_95_fu_1638;
reg   [7:0] tmp_V_96_fu_1642;
reg   [7:0] tmp_V_97_fu_1646;
reg   [7:0] tmp_V_98_fu_1650;
reg   [7:0] tmp_V_99_fu_1654;
reg   [7:0] tmp_V_100_fu_1658;
reg   [7:0] tmp_V_101_fu_1662;
reg   [7:0] tmp_V_102_fu_1666;
reg   [7:0] tmp_V_103_fu_1670;
reg   [7:0] tmp_V_104_fu_1674;
reg   [7:0] tmp_V_105_fu_1678;
reg   [7:0] tmp_V_106_fu_1682;
reg   [7:0] tmp_V_107_fu_1686;
reg   [7:0] tmp_V_108_fu_1690;
reg   [7:0] tmp_V_109_fu_1694;
reg   [7:0] tmp_V_110_fu_1698;
reg   [7:0] tmp_V_111_fu_1702;
reg   [7:0] tmp_V_112_fu_1706;
reg   [7:0] tmp_V_113_fu_1710;
reg   [7:0] tmp_V_114_fu_1714;
reg   [7:0] tmp_V_115_fu_1718;
reg   [7:0] tmp_V_116_fu_1722;
reg   [7:0] tmp_V_117_fu_1726;
reg   [7:0] tmp_V_118_fu_1730;
reg   [7:0] tmp_V_119_fu_1734;
reg   [7:0] tmp_V_120_fu_1738;
reg   [7:0] tmp_V_121_fu_1742;
reg   [7:0] tmp_V_122_fu_1746;
reg   [7:0] tmp_V_123_fu_1750;
reg   [7:0] tmp_V_124_fu_1754;
reg   [7:0] tmp_V_125_fu_1758;
reg   [7:0] tmp_V_126_fu_1762;
reg   [7:0] tmp_V_127_fu_1766;
reg   [7:0] tmp_V_128_fu_1770;
reg   [7:0] tmp_V_129_fu_1774;
reg   [7:0] tmp_V_130_fu_1778;
reg   [7:0] tmp_V_131_fu_1782;
reg   [7:0] tmp_V_132_fu_1786;
reg   [7:0] tmp_V_133_fu_1790;
reg   [7:0] tmp_V_134_fu_1794;
reg   [7:0] tmp_V_135_fu_1798;
reg   [7:0] tmp_V_136_fu_1802;
reg   [7:0] tmp_V_137_fu_1806;
reg   [7:0] tmp_V_138_fu_1810;
reg   [7:0] tmp_V_139_fu_1814;
reg   [7:0] tmp_V_140_fu_1818;
reg   [7:0] tmp_V_141_fu_1822;
reg   [7:0] tmp_V_142_fu_1826;
reg   [7:0] tmp_V_143_fu_1830;
reg   [7:0] tmp_V_144_fu_1834;
reg   [7:0] tmp_V_145_fu_1838;
reg   [7:0] tmp_V_146_fu_1842;
reg   [7:0] tmp_V_147_fu_1846;
reg   [7:0] tmp_V_148_fu_1850;
reg   [7:0] tmp_V_149_fu_1854;
reg   [7:0] tmp_V_150_fu_1858;
reg   [7:0] tmp_V_151_fu_1862;
reg   [7:0] tmp_V_152_fu_1866;
reg   [7:0] tmp_V_153_fu_1870;
reg   [7:0] tmp_V_154_fu_1874;
reg   [7:0] tmp_V_155_fu_1878;
reg   [7:0] tmp_V_156_fu_1882;
reg   [7:0] tmp_V_157_fu_1886;
reg   [7:0] tmp_V_158_fu_1890;
reg   [7:0] tmp_V_159_fu_1894;
reg   [7:0] tmp_V_160_fu_1898;
reg   [7:0] tmp_V_161_fu_1902;
reg   [7:0] tmp_V_162_fu_1906;
reg   [7:0] tmp_V_163_fu_1910;
reg   [7:0] tmp_V_164_fu_1914;
reg   [7:0] tmp_V_165_fu_1918;
reg   [7:0] tmp_V_166_fu_1922;
reg   [7:0] tmp_V_167_fu_1926;
reg   [7:0] tmp_V_168_fu_1930;
reg   [7:0] tmp_V_169_fu_1934;
reg   [7:0] tmp_V_170_fu_1938;
reg   [7:0] tmp_V_171_fu_1942;
reg   [7:0] tmp_V_172_fu_1946;
reg   [7:0] tmp_V_173_fu_1950;
reg   [7:0] tmp_V_174_fu_1954;
reg   [7:0] tmp_V_175_fu_1958;
reg   [7:0] tmp_V_176_fu_1962;
reg   [7:0] tmp_V_177_fu_1966;
reg   [7:0] tmp_V_178_fu_1970;
reg   [7:0] tmp_V_179_fu_1974;
reg   [7:0] tmp_V_180_fu_1978;
reg   [7:0] tmp_V_181_fu_1982;
reg   [7:0] tmp_V_182_fu_1986;
reg   [7:0] tmp_V_183_fu_1990;
reg   [7:0] tmp_V_184_fu_1994;
reg   [7:0] tmp_V_185_fu_1998;
reg   [7:0] tmp_V_186_fu_2002;
reg   [7:0] tmp_V_187_fu_2006;
reg   [7:0] tmp_V_188_fu_2010;
reg   [7:0] tmp_V_189_fu_2014;
reg   [7:0] tmp_V_190_fu_2018;
reg   [7:0] tmp_V_191_fu_2022;
reg   [7:0] tmp_V_192_fu_2026;
reg   [7:0] tmp_V_193_fu_2030;
reg   [7:0] tmp_V_194_fu_2034;
reg   [7:0] tmp_V_195_fu_2038;
reg   [7:0] tmp_V_196_fu_2042;
reg   [7:0] tmp_V_197_fu_2046;
reg   [7:0] tmp_V_198_fu_2050;
reg   [7:0] tmp_V_199_fu_2054;
reg   [7:0] tmp_V_200_fu_2058;
reg   [7:0] tmp_V_201_fu_2062;
reg   [7:0] tmp_V_202_fu_2066;
reg   [7:0] tmp_V_203_fu_2070;
reg   [7:0] tmp_V_204_fu_2074;
reg   [7:0] tmp_V_205_fu_2078;
reg   [7:0] tmp_V_206_fu_2082;
reg   [7:0] tmp_V_207_fu_2086;
reg   [7:0] tmp_V_208_fu_2090;
reg   [7:0] tmp_V_209_fu_2094;
reg   [7:0] tmp_V_210_fu_2098;
reg   [7:0] tmp_V_211_fu_2102;
reg   [7:0] tmp_V_212_fu_2106;
reg   [7:0] tmp_V_213_fu_2110;
reg   [7:0] tmp_V_214_fu_2114;
reg   [7:0] tmp_V_215_fu_2118;
reg   [7:0] tmp_V_216_fu_2122;
reg   [7:0] tmp_V_217_fu_2126;
reg   [7:0] tmp_V_218_fu_2130;
reg   [7:0] tmp_V_219_fu_2134;
reg   [7:0] tmp_V_220_fu_2138;
reg   [7:0] tmp_V_221_fu_2142;
reg   [7:0] tmp_V_222_fu_2146;
reg   [7:0] tmp_V_223_fu_2150;
reg   [7:0] tmp_V_224_fu_2154;
reg   [7:0] tmp_V_225_fu_2158;
reg   [7:0] tmp_V_226_fu_2162;
reg   [7:0] tmp_V_227_fu_2166;
reg   [7:0] tmp_V_228_fu_2170;
reg   [7:0] tmp_V_229_fu_2174;
reg   [7:0] tmp_V_230_fu_2178;
reg   [7:0] tmp_V_231_fu_2182;
reg   [7:0] tmp_V_232_fu_2186;
reg   [7:0] tmp_V_233_fu_2190;
reg   [7:0] tmp_V_234_fu_2194;
reg   [7:0] tmp_V_235_fu_2198;
reg   [7:0] tmp_V_236_fu_2202;
reg   [7:0] tmp_V_237_fu_2206;
reg   [7:0] tmp_V_238_fu_2210;
reg   [7:0] tmp_V_239_fu_2214;
reg   [7:0] tmp_V_240_fu_2218;
reg   [7:0] tmp_V_241_fu_2222;
reg   [7:0] tmp_V_242_fu_2226;
reg   [7:0] tmp_V_243_fu_2230;
reg   [7:0] tmp_V_244_fu_2234;
reg   [7:0] tmp_V_245_fu_2238;
reg   [7:0] tmp_V_246_fu_2242;
reg   [7:0] tmp_V_247_fu_2246;
reg   [7:0] tmp_V_248_fu_2250;
reg   [7:0] tmp_V_249_fu_2254;
reg   [7:0] tmp_V_250_fu_2258;
reg   [7:0] tmp_V_251_fu_2262;
reg   [7:0] tmp_V_252_fu_2266;
reg   [7:0] tmp_V_253_fu_2270;
reg   [7:0] tmp_V_254_fu_2274;
reg   [7:0] tmp_V_255_fu_2278;
reg   [7:0] tmp_V_256_fu_2282;
reg   [7:0] tmp_V_257_fu_2286;
reg   [7:0] tmp_V_258_fu_2290;
reg   [7:0] tmp_V_259_fu_2294;
reg   [7:0] tmp_V_260_fu_2298;
reg   [7:0] tmp_V_261_fu_2302;
reg   [7:0] tmp_V_262_fu_2306;
reg   [7:0] tmp_V_263_fu_2310;
reg   [7:0] tmp_V_264_fu_2314;
reg   [7:0] tmp_V_265_fu_2318;
reg   [7:0] tmp_V_266_fu_2322;
reg   [7:0] tmp_V_267_fu_2326;
reg   [7:0] tmp_V_268_fu_2330;
reg   [7:0] tmp_V_269_fu_2334;
reg   [7:0] tmp_V_270_fu_2338;
reg   [7:0] tmp_V_271_fu_2342;
reg   [7:0] tmp_V_272_fu_2346;
reg   [7:0] tmp_V_273_fu_2350;
reg   [7:0] tmp_V_274_fu_2354;
reg   [7:0] tmp_V_275_fu_2358;
reg   [7:0] tmp_V_276_fu_2362;
reg   [7:0] tmp_V_277_fu_2366;
reg   [7:0] tmp_V_278_fu_2370;
reg   [7:0] tmp_V_279_fu_2374;
reg   [7:0] tmp_V_280_fu_2378;
reg   [7:0] tmp_V_281_fu_2382;
reg   [7:0] tmp_V_282_fu_2386;
reg   [7:0] tmp_V_283_fu_2390;
reg   [7:0] tmp_V_284_fu_2394;
reg   [7:0] tmp_V_285_fu_2398;
reg   [7:0] tmp_V_286_fu_2402;
reg   [7:0] tmp_V_287_fu_2406;
reg   [7:0] tmp_V_288_fu_2410;
reg   [7:0] tmp_V_289_fu_2414;
reg   [7:0] tmp_V_290_fu_2418;
reg   [7:0] tmp_V_291_fu_2422;
reg   [7:0] tmp_V_292_fu_2426;
reg   [7:0] tmp_V_293_fu_2430;
reg   [7:0] tmp_V_294_fu_2434;
reg   [7:0] tmp_V_295_fu_2438;
reg   [7:0] tmp_V_296_fu_2442;
reg   [7:0] tmp_V_297_fu_2446;
reg   [7:0] tmp_V_298_fu_2450;
reg   [7:0] tmp_V_299_fu_2454;
reg   [7:0] tmp_V_300_fu_2458;
reg   [7:0] tmp_V_301_fu_2462;
reg   [7:0] tmp_V_302_fu_2466;
reg   [7:0] tmp_V_303_fu_2470;
reg   [7:0] tmp_V_304_fu_2474;
reg   [7:0] tmp_V_305_fu_2478;
reg   [7:0] tmp_V_306_fu_2482;
reg   [7:0] tmp_V_307_fu_2486;
reg   [7:0] tmp_V_308_fu_2490;
reg   [7:0] tmp_V_309_fu_2494;
reg   [7:0] tmp_V_310_fu_2498;
reg   [7:0] tmp_V_311_fu_2502;
reg   [7:0] tmp_V_312_fu_2506;
reg   [7:0] tmp_V_313_fu_2510;
reg   [7:0] tmp_V_314_fu_2514;
reg   [7:0] tmp_V_315_fu_2518;
reg   [7:0] tmp_V_316_fu_2522;
reg   [7:0] tmp_V_317_fu_2526;
reg   [7:0] tmp_V_318_fu_2530;
reg   [7:0] tmp_V_319_fu_2534;
reg   [7:0] tmp_V_320_fu_2538;
reg   [7:0] tmp_V_321_fu_2542;
reg   [7:0] tmp_V_322_fu_2546;
reg   [7:0] tmp_V_323_fu_2550;
reg   [7:0] tmp_V_324_fu_2554;
reg   [7:0] tmp_V_325_fu_2558;
reg   [7:0] tmp_V_326_fu_2562;
reg   [7:0] tmp_V_327_fu_2566;
reg   [7:0] tmp_V_328_fu_2570;
reg   [7:0] tmp_V_329_fu_2574;
reg   [7:0] tmp_V_330_fu_2578;
reg   [7:0] tmp_V_331_fu_2582;
reg   [7:0] tmp_V_332_fu_2586;
reg   [7:0] tmp_V_333_fu_2590;
reg   [7:0] tmp_V_334_fu_2594;
reg   [7:0] tmp_V_335_fu_2598;
reg   [7:0] tmp_V_336_fu_2602;
reg   [7:0] tmp_V_337_fu_2606;
reg   [7:0] tmp_V_338_fu_2610;
reg   [7:0] tmp_V_339_fu_2614;
reg   [7:0] tmp_V_340_fu_2618;
reg   [7:0] tmp_V_341_fu_2622;
reg   [7:0] tmp_V_342_fu_2626;
reg   [7:0] tmp_V_343_fu_2630;
reg   [7:0] tmp_V_344_fu_2634;
reg   [7:0] tmp_V_345_fu_2638;
reg   [7:0] tmp_V_346_fu_2642;
reg   [7:0] tmp_V_347_fu_2646;
reg   [7:0] tmp_V_348_fu_2650;
reg   [7:0] tmp_V_349_fu_2654;
reg   [7:0] tmp_V_350_fu_2658;
reg   [7:0] tmp_V_351_fu_2662;
reg   [7:0] tmp_V_352_fu_2666;
reg   [7:0] tmp_V_353_fu_2670;
reg   [7:0] tmp_V_354_fu_2674;
reg   [7:0] tmp_V_355_fu_2678;
reg   [7:0] tmp_V_356_fu_2682;
reg   [7:0] tmp_V_357_fu_2686;
reg   [7:0] tmp_V_358_fu_2690;
reg   [7:0] tmp_V_359_fu_2694;
reg   [7:0] tmp_V_360_fu_2698;
reg   [7:0] tmp_V_361_fu_2702;
reg   [7:0] tmp_V_362_fu_2706;
reg   [7:0] tmp_V_363_fu_2710;
reg   [7:0] tmp_V_364_fu_2714;
reg   [7:0] tmp_V_365_fu_2718;
reg   [7:0] tmp_V_366_fu_2722;
reg   [7:0] tmp_V_367_fu_2726;
reg   [7:0] tmp_V_368_fu_2730;
reg   [7:0] tmp_V_369_fu_2734;
reg   [7:0] tmp_V_370_fu_2738;
reg   [7:0] tmp_V_371_fu_2742;
reg   [7:0] tmp_V_372_fu_2746;
reg   [7:0] tmp_V_373_fu_2750;
reg   [7:0] tmp_V_374_fu_2754;
reg   [7:0] tmp_V_375_fu_2758;
reg   [7:0] tmp_V_376_fu_2762;
reg   [7:0] tmp_V_377_fu_2766;
reg   [7:0] tmp_V_378_fu_2770;
reg   [7:0] tmp_V_379_fu_2774;
reg   [7:0] tmp_V_380_fu_2778;
reg   [7:0] tmp_V_381_fu_2782;
reg   [7:0] tmp_V_382_fu_2786;
reg   [7:0] tmp_V_383_fu_2790;
reg   [7:0] tmp_V_384_fu_2794;
reg   [7:0] tmp_V_385_fu_2798;
reg   [7:0] tmp_V_386_fu_2802;
reg   [7:0] tmp_V_387_fu_2806;
reg   [7:0] tmp_V_388_fu_2810;
reg   [7:0] tmp_V_389_fu_2814;
reg   [7:0] tmp_V_390_fu_2818;
reg   [7:0] tmp_V_391_fu_2822;
reg   [7:0] tmp_V_392_fu_2826;
reg   [7:0] tmp_V_393_fu_2830;
reg   [7:0] tmp_V_394_fu_2834;
reg   [7:0] tmp_V_395_fu_2838;
reg   [7:0] tmp_V_396_fu_2842;
reg   [7:0] tmp_V_397_fu_2846;
reg   [7:0] tmp_V_398_fu_2850;
reg   [7:0] tmp_V_399_fu_2854;
reg   [7:0] tmp_V_400_fu_2858;
reg   [7:0] tmp_V_401_fu_2862;
reg   [7:0] tmp_V_402_fu_2866;
reg   [7:0] tmp_V_403_fu_2870;
reg   [7:0] tmp_V_404_fu_2874;
reg   [7:0] tmp_V_405_fu_2878;
reg   [7:0] tmp_V_406_fu_2882;
reg   [7:0] tmp_V_407_fu_2886;
reg   [7:0] tmp_V_408_fu_2890;
reg   [7:0] tmp_V_409_fu_2894;
reg   [7:0] tmp_V_410_fu_2898;
reg   [7:0] tmp_V_411_fu_2902;
reg   [7:0] tmp_V_412_fu_2906;
reg   [7:0] tmp_V_413_fu_2910;
reg   [7:0] tmp_V_414_fu_2914;
reg   [7:0] tmp_V_415_fu_2918;
reg   [7:0] tmp_V_416_fu_2922;
reg   [7:0] tmp_V_417_fu_2926;
reg   [7:0] tmp_V_418_fu_2930;
reg   [7:0] tmp_V_419_fu_2934;
reg   [7:0] tmp_V_420_fu_2938;
reg   [7:0] tmp_V_421_fu_2942;
reg   [7:0] tmp_V_422_fu_2946;
reg   [7:0] tmp_V_423_fu_2950;
reg   [7:0] tmp_V_424_fu_2954;
reg   [7:0] tmp_V_425_fu_2958;
reg   [7:0] tmp_V_426_fu_2962;
reg   [7:0] tmp_V_427_fu_2966;
reg   [7:0] tmp_V_428_fu_2970;
reg   [7:0] tmp_V_429_fu_2974;
reg   [7:0] tmp_V_430_fu_2978;
reg   [7:0] tmp_V_431_fu_2982;
reg   [7:0] tmp_V_432_fu_2986;
reg   [7:0] tmp_V_433_fu_2990;
reg   [7:0] tmp_V_434_fu_2994;
reg   [7:0] tmp_V_435_fu_2998;
reg   [7:0] tmp_V_436_fu_3002;
reg   [7:0] tmp_V_437_fu_3006;
reg   [7:0] tmp_V_438_fu_3010;
reg   [7:0] tmp_V_439_fu_3014;
reg   [7:0] tmp_V_440_fu_3018;
reg   [7:0] tmp_V_441_fu_3022;
reg   [7:0] tmp_V_442_fu_3026;
reg   [7:0] tmp_V_443_fu_3030;
reg   [7:0] tmp_V_444_fu_3034;
reg   [7:0] tmp_V_445_fu_3038;
reg   [7:0] tmp_V_446_fu_3042;
reg   [7:0] tmp_V_447_fu_3046;
reg   [7:0] tmp_V_448_fu_3050;
reg   [7:0] tmp_V_449_fu_3054;
reg   [7:0] tmp_V_450_fu_3058;
reg   [7:0] tmp_V_451_fu_3062;
reg   [7:0] tmp_V_452_fu_3066;
reg   [7:0] tmp_V_453_fu_3070;
reg   [7:0] tmp_V_454_fu_3074;
reg   [7:0] tmp_V_455_fu_3078;
reg   [7:0] tmp_V_456_fu_3082;
reg   [7:0] tmp_V_457_fu_3086;
reg   [7:0] tmp_V_458_fu_3090;
reg   [7:0] tmp_V_459_fu_3094;
reg   [7:0] tmp_V_460_fu_3098;
reg   [7:0] tmp_V_461_fu_3102;
reg   [7:0] tmp_V_462_fu_3106;
reg   [7:0] tmp_V_463_fu_3110;
reg   [7:0] tmp_V_464_fu_3114;
reg   [7:0] tmp_V_465_fu_3118;
reg   [7:0] tmp_V_466_fu_3122;
reg   [7:0] tmp_V_467_fu_3126;
reg   [7:0] tmp_V_468_fu_3130;
reg   [7:0] tmp_V_469_fu_3134;
reg   [7:0] tmp_V_470_fu_3138;
reg   [7:0] tmp_V_471_fu_3142;
reg   [7:0] tmp_V_472_fu_3146;
reg   [7:0] tmp_V_473_fu_3150;
reg   [7:0] tmp_V_474_fu_3154;
reg   [7:0] tmp_V_475_fu_3158;
reg   [7:0] tmp_V_476_fu_3162;
reg   [7:0] tmp_V_477_fu_3166;
reg   [7:0] tmp_V_478_fu_3170;
reg   [7:0] tmp_V_479_fu_3174;
reg   [7:0] tmp_V_480_fu_3178;
reg   [7:0] tmp_V_481_fu_3182;
reg   [7:0] tmp_V_482_fu_3186;
reg   [7:0] tmp_V_483_fu_3190;
reg   [7:0] tmp_V_484_fu_3194;
reg   [7:0] tmp_V_485_fu_3198;
reg   [7:0] tmp_V_486_fu_3202;
reg   [7:0] tmp_V_487_fu_3206;
reg   [7:0] tmp_V_488_fu_3210;
reg   [7:0] tmp_V_489_fu_3214;
reg   [7:0] tmp_V_490_fu_3218;
reg   [7:0] tmp_V_491_fu_3222;
reg   [7:0] tmp_V_492_fu_3226;
reg   [7:0] tmp_V_493_fu_3230;
reg   [7:0] tmp_V_494_fu_3234;
reg   [7:0] tmp_V_495_fu_3238;
reg   [7:0] tmp_V_496_fu_3242;
reg   [7:0] tmp_V_497_fu_3246;
reg   [7:0] tmp_V_498_fu_3250;
reg   [7:0] tmp_V_499_fu_3254;
reg   [7:0] tmp_V_500_fu_3258;
reg   [7:0] tmp_V_501_fu_3262;
reg   [7:0] tmp_V_502_fu_3266;
reg   [7:0] tmp_V_503_fu_3270;
reg   [7:0] tmp_V_504_fu_3274;
reg   [7:0] tmp_V_505_fu_3278;
reg   [7:0] tmp_V_506_fu_3282;
reg   [7:0] tmp_V_507_fu_3286;
reg   [7:0] tmp_V_508_fu_3290;
reg   [7:0] tmp_V_509_fu_3294;
reg   [7:0] tmp_V_510_fu_3298;
reg   [7:0] tmp_V_511_fu_3302;
reg   [7:0] tmp_V_512_fu_3306;
reg   [7:0] tmp_V_513_fu_3310;
reg   [7:0] tmp_V_514_fu_3314;
reg   [7:0] tmp_V_515_fu_3318;
reg   [7:0] tmp_V_516_fu_3322;
reg   [7:0] tmp_V_517_fu_3326;
reg   [7:0] tmp_V_518_fu_3330;
reg   [7:0] tmp_V_519_fu_3334;
reg   [7:0] tmp_V_520_fu_3338;
reg   [7:0] tmp_V_521_fu_3342;
reg   [7:0] tmp_V_522_fu_3346;
reg   [7:0] tmp_V_523_fu_3350;
reg   [7:0] tmp_V_524_fu_3354;
reg   [7:0] tmp_V_525_fu_3358;
reg   [7:0] tmp_V_526_fu_3362;
reg   [7:0] tmp_V_527_fu_3366;
reg   [7:0] tmp_V_528_fu_3370;
reg   [7:0] tmp_V_529_fu_3374;
reg   [7:0] tmp_V_530_fu_3378;
reg   [7:0] tmp_V_531_fu_3382;
reg   [7:0] tmp_V_532_fu_3386;
reg   [7:0] tmp_V_533_fu_3390;
reg   [7:0] tmp_V_534_fu_3394;
reg   [7:0] tmp_V_535_fu_3398;
reg   [7:0] tmp_V_536_fu_3402;
reg   [7:0] tmp_V_537_fu_3406;
reg   [7:0] tmp_V_538_fu_3410;
reg   [7:0] tmp_V_539_fu_3414;
reg   [7:0] tmp_V_540_fu_3418;
reg   [7:0] tmp_V_541_fu_3422;
reg   [7:0] tmp_V_542_fu_3426;
reg   [7:0] tmp_V_543_fu_3430;
reg   [7:0] tmp_V_544_fu_3434;
reg   [7:0] tmp_V_545_fu_3438;
reg   [7:0] tmp_V_546_fu_3442;
reg   [7:0] tmp_V_547_fu_3446;
reg   [7:0] tmp_V_548_fu_3450;
reg   [7:0] tmp_V_549_fu_3454;
reg   [7:0] tmp_V_550_fu_3458;
reg   [7:0] tmp_V_551_fu_3462;
reg   [7:0] tmp_V_552_fu_3466;
reg   [7:0] tmp_V_553_fu_3470;
reg   [7:0] tmp_V_554_fu_3474;
reg   [7:0] tmp_V_555_fu_3478;
reg   [7:0] tmp_V_556_fu_3482;
reg   [7:0] tmp_V_557_fu_3486;
reg   [7:0] tmp_V_558_fu_3490;
reg   [7:0] tmp_V_559_fu_3494;
reg   [7:0] tmp_V_560_fu_3498;
reg   [7:0] tmp_V_561_fu_3502;
reg   [7:0] tmp_V_562_fu_3506;
reg   [7:0] tmp_V_563_fu_3510;
reg   [7:0] tmp_V_564_fu_3514;
reg   [7:0] tmp_V_565_fu_3518;
reg   [7:0] tmp_V_566_fu_3522;
reg   [7:0] tmp_V_567_fu_3526;
reg   [7:0] tmp_V_568_fu_3530;
reg   [7:0] tmp_V_569_fu_3534;
reg   [7:0] tmp_V_570_fu_3538;
reg   [7:0] tmp_V_571_fu_3542;
reg   [7:0] tmp_V_572_fu_3546;
reg   [7:0] tmp_V_573_fu_3550;
reg   [7:0] tmp_V_574_fu_3554;
reg   [7:0] tmp_V_575_fu_3558;
reg   [7:0] tmp_V_576_fu_3562;
reg   [31:0] nf_0_fu_3566;
wire   [31:0] select_ln301_fu_10945_p3;
reg   [31:0] ap_sig_allocacmp_nf_0_load_1;
reg    ap_block_pp0_stage0_01001;
wire   [9:0] inElem_V_1_fu_6525_p577;
wire   [3:0] trunc_ln647_1_fu_10707_p1;
wire  signed [3:0] mul_ln1352_fu_10718_p0;
wire  signed [7:0] sext_ln215_1_fu_10714_p1;
wire  signed [7:0] mul_ln1352_fu_10718_p2;
wire   [3:0] arg_V_read_assign_1_fu_10728_p4;
wire  signed [3:0] mul_ln1352_1_fu_10745_p0;
wire  signed [7:0] sext_ln215_3_fu_10741_p1;
wire  signed [7:0] mul_ln1352_1_fu_10745_p2;
wire  signed [8:0] sext_ln700_fu_10751_p1;
wire  signed [8:0] sext_ln170_fu_10724_p1;
wire   [8:0] add_ln700_fu_10755_p2;
wire   [23:0] select_ln271_3_fu_10700_p3;
wire  signed [23:0] sext_ln700_1_fu_10761_p1;
wire  signed [3:0] mul_ln1352_2_fu_10774_p0;
wire  signed [7:0] mul_ln1352_2_fu_10774_p2;
wire  signed [3:0] mul_ln1352_3_fu_10787_p0;
wire  signed [7:0] mul_ln1352_3_fu_10787_p2;
wire  signed [8:0] sext_ln700_2_fu_10793_p1;
wire  signed [8:0] sext_ln170_1_fu_10780_p1;
wire   [8:0] add_ln700_2_fu_10797_p2;
wire   [23:0] select_ln271_2_fu_10693_p3;
wire  signed [23:0] sext_ln700_3_fu_10803_p1;
wire  signed [3:0] mul_ln1352_4_fu_10816_p0;
wire  signed [7:0] mul_ln1352_4_fu_10816_p2;
wire  signed [3:0] mul_ln1352_5_fu_10829_p0;
wire  signed [7:0] mul_ln1352_5_fu_10829_p2;
wire  signed [8:0] sext_ln700_4_fu_10835_p1;
wire  signed [8:0] sext_ln170_2_fu_10822_p1;
wire   [8:0] add_ln700_4_fu_10839_p2;
wire   [23:0] select_ln271_1_fu_10686_p3;
wire  signed [23:0] sext_ln700_5_fu_10845_p1;
wire  signed [3:0] mul_ln1352_6_fu_10858_p0;
wire  signed [7:0] mul_ln1352_6_fu_10858_p2;
wire  signed [3:0] mul_ln1352_7_fu_10871_p0;
wire  signed [7:0] mul_ln1352_7_fu_10871_p2;
wire  signed [8:0] sext_ln700_6_fu_10877_p1;
wire  signed [8:0] sext_ln170_3_fu_10864_p1;
wire   [8:0] add_ln700_6_fu_10881_p2;
wire   [23:0] select_ln271_fu_10679_p3;
wire  signed [23:0] sext_ln700_7_fu_10887_p1;
wire   [31:0] nf_fu_10933_p2;
wire   [0:0] icmp_ln301_fu_10939_p2;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

StreamingFCLayer_Batch_0_StreamingFCLayer_bkb #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 8 ),
    .din2_WIDTH( 8 ),
    .din3_WIDTH( 8 ),
    .din4_WIDTH( 8 ),
    .din5_WIDTH( 8 ),
    .din6_WIDTH( 8 ),
    .din7_WIDTH( 8 ),
    .din8_WIDTH( 8 ),
    .din9_WIDTH( 8 ),
    .din10_WIDTH( 8 ),
    .din11_WIDTH( 8 ),
    .din12_WIDTH( 8 ),
    .din13_WIDTH( 8 ),
    .din14_WIDTH( 8 ),
    .din15_WIDTH( 8 ),
    .din16_WIDTH( 8 ),
    .din17_WIDTH( 8 ),
    .din18_WIDTH( 8 ),
    .din19_WIDTH( 8 ),
    .din20_WIDTH( 8 ),
    .din21_WIDTH( 8 ),
    .din22_WIDTH( 8 ),
    .din23_WIDTH( 8 ),
    .din24_WIDTH( 8 ),
    .din25_WIDTH( 8 ),
    .din26_WIDTH( 8 ),
    .din27_WIDTH( 8 ),
    .din28_WIDTH( 8 ),
    .din29_WIDTH( 8 ),
    .din30_WIDTH( 8 ),
    .din31_WIDTH( 8 ),
    .din32_WIDTH( 8 ),
    .din33_WIDTH( 8 ),
    .din34_WIDTH( 8 ),
    .din35_WIDTH( 8 ),
    .din36_WIDTH( 8 ),
    .din37_WIDTH( 8 ),
    .din38_WIDTH( 8 ),
    .din39_WIDTH( 8 ),
    .din40_WIDTH( 8 ),
    .din41_WIDTH( 8 ),
    .din42_WIDTH( 8 ),
    .din43_WIDTH( 8 ),
    .din44_WIDTH( 8 ),
    .din45_WIDTH( 8 ),
    .din46_WIDTH( 8 ),
    .din47_WIDTH( 8 ),
    .din48_WIDTH( 8 ),
    .din49_WIDTH( 8 ),
    .din50_WIDTH( 8 ),
    .din51_WIDTH( 8 ),
    .din52_WIDTH( 8 ),
    .din53_WIDTH( 8 ),
    .din54_WIDTH( 8 ),
    .din55_WIDTH( 8 ),
    .din56_WIDTH( 8 ),
    .din57_WIDTH( 8 ),
    .din58_WIDTH( 8 ),
    .din59_WIDTH( 8 ),
    .din60_WIDTH( 8 ),
    .din61_WIDTH( 8 ),
    .din62_WIDTH( 8 ),
    .din63_WIDTH( 8 ),
    .din64_WIDTH( 8 ),
    .din65_WIDTH( 8 ),
    .din66_WIDTH( 8 ),
    .din67_WIDTH( 8 ),
    .din68_WIDTH( 8 ),
    .din69_WIDTH( 8 ),
    .din70_WIDTH( 8 ),
    .din71_WIDTH( 8 ),
    .din72_WIDTH( 8 ),
    .din73_WIDTH( 8 ),
    .din74_WIDTH( 8 ),
    .din75_WIDTH( 8 ),
    .din76_WIDTH( 8 ),
    .din77_WIDTH( 8 ),
    .din78_WIDTH( 8 ),
    .din79_WIDTH( 8 ),
    .din80_WIDTH( 8 ),
    .din81_WIDTH( 8 ),
    .din82_WIDTH( 8 ),
    .din83_WIDTH( 8 ),
    .din84_WIDTH( 8 ),
    .din85_WIDTH( 8 ),
    .din86_WIDTH( 8 ),
    .din87_WIDTH( 8 ),
    .din88_WIDTH( 8 ),
    .din89_WIDTH( 8 ),
    .din90_WIDTH( 8 ),
    .din91_WIDTH( 8 ),
    .din92_WIDTH( 8 ),
    .din93_WIDTH( 8 ),
    .din94_WIDTH( 8 ),
    .din95_WIDTH( 8 ),
    .din96_WIDTH( 8 ),
    .din97_WIDTH( 8 ),
    .din98_WIDTH( 8 ),
    .din99_WIDTH( 8 ),
    .din100_WIDTH( 8 ),
    .din101_WIDTH( 8 ),
    .din102_WIDTH( 8 ),
    .din103_WIDTH( 8 ),
    .din104_WIDTH( 8 ),
    .din105_WIDTH( 8 ),
    .din106_WIDTH( 8 ),
    .din107_WIDTH( 8 ),
    .din108_WIDTH( 8 ),
    .din109_WIDTH( 8 ),
    .din110_WIDTH( 8 ),
    .din111_WIDTH( 8 ),
    .din112_WIDTH( 8 ),
    .din113_WIDTH( 8 ),
    .din114_WIDTH( 8 ),
    .din115_WIDTH( 8 ),
    .din116_WIDTH( 8 ),
    .din117_WIDTH( 8 ),
    .din118_WIDTH( 8 ),
    .din119_WIDTH( 8 ),
    .din120_WIDTH( 8 ),
    .din121_WIDTH( 8 ),
    .din122_WIDTH( 8 ),
    .din123_WIDTH( 8 ),
    .din124_WIDTH( 8 ),
    .din125_WIDTH( 8 ),
    .din126_WIDTH( 8 ),
    .din127_WIDTH( 8 ),
    .din128_WIDTH( 8 ),
    .din129_WIDTH( 8 ),
    .din130_WIDTH( 8 ),
    .din131_WIDTH( 8 ),
    .din132_WIDTH( 8 ),
    .din133_WIDTH( 8 ),
    .din134_WIDTH( 8 ),
    .din135_WIDTH( 8 ),
    .din136_WIDTH( 8 ),
    .din137_WIDTH( 8 ),
    .din138_WIDTH( 8 ),
    .din139_WIDTH( 8 ),
    .din140_WIDTH( 8 ),
    .din141_WIDTH( 8 ),
    .din142_WIDTH( 8 ),
    .din143_WIDTH( 8 ),
    .din144_WIDTH( 8 ),
    .din145_WIDTH( 8 ),
    .din146_WIDTH( 8 ),
    .din147_WIDTH( 8 ),
    .din148_WIDTH( 8 ),
    .din149_WIDTH( 8 ),
    .din150_WIDTH( 8 ),
    .din151_WIDTH( 8 ),
    .din152_WIDTH( 8 ),
    .din153_WIDTH( 8 ),
    .din154_WIDTH( 8 ),
    .din155_WIDTH( 8 ),
    .din156_WIDTH( 8 ),
    .din157_WIDTH( 8 ),
    .din158_WIDTH( 8 ),
    .din159_WIDTH( 8 ),
    .din160_WIDTH( 8 ),
    .din161_WIDTH( 8 ),
    .din162_WIDTH( 8 ),
    .din163_WIDTH( 8 ),
    .din164_WIDTH( 8 ),
    .din165_WIDTH( 8 ),
    .din166_WIDTH( 8 ),
    .din167_WIDTH( 8 ),
    .din168_WIDTH( 8 ),
    .din169_WIDTH( 8 ),
    .din170_WIDTH( 8 ),
    .din171_WIDTH( 8 ),
    .din172_WIDTH( 8 ),
    .din173_WIDTH( 8 ),
    .din174_WIDTH( 8 ),
    .din175_WIDTH( 8 ),
    .din176_WIDTH( 8 ),
    .din177_WIDTH( 8 ),
    .din178_WIDTH( 8 ),
    .din179_WIDTH( 8 ),
    .din180_WIDTH( 8 ),
    .din181_WIDTH( 8 ),
    .din182_WIDTH( 8 ),
    .din183_WIDTH( 8 ),
    .din184_WIDTH( 8 ),
    .din185_WIDTH( 8 ),
    .din186_WIDTH( 8 ),
    .din187_WIDTH( 8 ),
    .din188_WIDTH( 8 ),
    .din189_WIDTH( 8 ),
    .din190_WIDTH( 8 ),
    .din191_WIDTH( 8 ),
    .din192_WIDTH( 8 ),
    .din193_WIDTH( 8 ),
    .din194_WIDTH( 8 ),
    .din195_WIDTH( 8 ),
    .din196_WIDTH( 8 ),
    .din197_WIDTH( 8 ),
    .din198_WIDTH( 8 ),
    .din199_WIDTH( 8 ),
    .din200_WIDTH( 8 ),
    .din201_WIDTH( 8 ),
    .din202_WIDTH( 8 ),
    .din203_WIDTH( 8 ),
    .din204_WIDTH( 8 ),
    .din205_WIDTH( 8 ),
    .din206_WIDTH( 8 ),
    .din207_WIDTH( 8 ),
    .din208_WIDTH( 8 ),
    .din209_WIDTH( 8 ),
    .din210_WIDTH( 8 ),
    .din211_WIDTH( 8 ),
    .din212_WIDTH( 8 ),
    .din213_WIDTH( 8 ),
    .din214_WIDTH( 8 ),
    .din215_WIDTH( 8 ),
    .din216_WIDTH( 8 ),
    .din217_WIDTH( 8 ),
    .din218_WIDTH( 8 ),
    .din219_WIDTH( 8 ),
    .din220_WIDTH( 8 ),
    .din221_WIDTH( 8 ),
    .din222_WIDTH( 8 ),
    .din223_WIDTH( 8 ),
    .din224_WIDTH( 8 ),
    .din225_WIDTH( 8 ),
    .din226_WIDTH( 8 ),
    .din227_WIDTH( 8 ),
    .din228_WIDTH( 8 ),
    .din229_WIDTH( 8 ),
    .din230_WIDTH( 8 ),
    .din231_WIDTH( 8 ),
    .din232_WIDTH( 8 ),
    .din233_WIDTH( 8 ),
    .din234_WIDTH( 8 ),
    .din235_WIDTH( 8 ),
    .din236_WIDTH( 8 ),
    .din237_WIDTH( 8 ),
    .din238_WIDTH( 8 ),
    .din239_WIDTH( 8 ),
    .din240_WIDTH( 8 ),
    .din241_WIDTH( 8 ),
    .din242_WIDTH( 8 ),
    .din243_WIDTH( 8 ),
    .din244_WIDTH( 8 ),
    .din245_WIDTH( 8 ),
    .din246_WIDTH( 8 ),
    .din247_WIDTH( 8 ),
    .din248_WIDTH( 8 ),
    .din249_WIDTH( 8 ),
    .din250_WIDTH( 8 ),
    .din251_WIDTH( 8 ),
    .din252_WIDTH( 8 ),
    .din253_WIDTH( 8 ),
    .din254_WIDTH( 8 ),
    .din255_WIDTH( 8 ),
    .din256_WIDTH( 8 ),
    .din257_WIDTH( 8 ),
    .din258_WIDTH( 8 ),
    .din259_WIDTH( 8 ),
    .din260_WIDTH( 8 ),
    .din261_WIDTH( 8 ),
    .din262_WIDTH( 8 ),
    .din263_WIDTH( 8 ),
    .din264_WIDTH( 8 ),
    .din265_WIDTH( 8 ),
    .din266_WIDTH( 8 ),
    .din267_WIDTH( 8 ),
    .din268_WIDTH( 8 ),
    .din269_WIDTH( 8 ),
    .din270_WIDTH( 8 ),
    .din271_WIDTH( 8 ),
    .din272_WIDTH( 8 ),
    .din273_WIDTH( 8 ),
    .din274_WIDTH( 8 ),
    .din275_WIDTH( 8 ),
    .din276_WIDTH( 8 ),
    .din277_WIDTH( 8 ),
    .din278_WIDTH( 8 ),
    .din279_WIDTH( 8 ),
    .din280_WIDTH( 8 ),
    .din281_WIDTH( 8 ),
    .din282_WIDTH( 8 ),
    .din283_WIDTH( 8 ),
    .din284_WIDTH( 8 ),
    .din285_WIDTH( 8 ),
    .din286_WIDTH( 8 ),
    .din287_WIDTH( 8 ),
    .din288_WIDTH( 8 ),
    .din289_WIDTH( 8 ),
    .din290_WIDTH( 8 ),
    .din291_WIDTH( 8 ),
    .din292_WIDTH( 8 ),
    .din293_WIDTH( 8 ),
    .din294_WIDTH( 8 ),
    .din295_WIDTH( 8 ),
    .din296_WIDTH( 8 ),
    .din297_WIDTH( 8 ),
    .din298_WIDTH( 8 ),
    .din299_WIDTH( 8 ),
    .din300_WIDTH( 8 ),
    .din301_WIDTH( 8 ),
    .din302_WIDTH( 8 ),
    .din303_WIDTH( 8 ),
    .din304_WIDTH( 8 ),
    .din305_WIDTH( 8 ),
    .din306_WIDTH( 8 ),
    .din307_WIDTH( 8 ),
    .din308_WIDTH( 8 ),
    .din309_WIDTH( 8 ),
    .din310_WIDTH( 8 ),
    .din311_WIDTH( 8 ),
    .din312_WIDTH( 8 ),
    .din313_WIDTH( 8 ),
    .din314_WIDTH( 8 ),
    .din315_WIDTH( 8 ),
    .din316_WIDTH( 8 ),
    .din317_WIDTH( 8 ),
    .din318_WIDTH( 8 ),
    .din319_WIDTH( 8 ),
    .din320_WIDTH( 8 ),
    .din321_WIDTH( 8 ),
    .din322_WIDTH( 8 ),
    .din323_WIDTH( 8 ),
    .din324_WIDTH( 8 ),
    .din325_WIDTH( 8 ),
    .din326_WIDTH( 8 ),
    .din327_WIDTH( 8 ),
    .din328_WIDTH( 8 ),
    .din329_WIDTH( 8 ),
    .din330_WIDTH( 8 ),
    .din331_WIDTH( 8 ),
    .din332_WIDTH( 8 ),
    .din333_WIDTH( 8 ),
    .din334_WIDTH( 8 ),
    .din335_WIDTH( 8 ),
    .din336_WIDTH( 8 ),
    .din337_WIDTH( 8 ),
    .din338_WIDTH( 8 ),
    .din339_WIDTH( 8 ),
    .din340_WIDTH( 8 ),
    .din341_WIDTH( 8 ),
    .din342_WIDTH( 8 ),
    .din343_WIDTH( 8 ),
    .din344_WIDTH( 8 ),
    .din345_WIDTH( 8 ),
    .din346_WIDTH( 8 ),
    .din347_WIDTH( 8 ),
    .din348_WIDTH( 8 ),
    .din349_WIDTH( 8 ),
    .din350_WIDTH( 8 ),
    .din351_WIDTH( 8 ),
    .din352_WIDTH( 8 ),
    .din353_WIDTH( 8 ),
    .din354_WIDTH( 8 ),
    .din355_WIDTH( 8 ),
    .din356_WIDTH( 8 ),
    .din357_WIDTH( 8 ),
    .din358_WIDTH( 8 ),
    .din359_WIDTH( 8 ),
    .din360_WIDTH( 8 ),
    .din361_WIDTH( 8 ),
    .din362_WIDTH( 8 ),
    .din363_WIDTH( 8 ),
    .din364_WIDTH( 8 ),
    .din365_WIDTH( 8 ),
    .din366_WIDTH( 8 ),
    .din367_WIDTH( 8 ),
    .din368_WIDTH( 8 ),
    .din369_WIDTH( 8 ),
    .din370_WIDTH( 8 ),
    .din371_WIDTH( 8 ),
    .din372_WIDTH( 8 ),
    .din373_WIDTH( 8 ),
    .din374_WIDTH( 8 ),
    .din375_WIDTH( 8 ),
    .din376_WIDTH( 8 ),
    .din377_WIDTH( 8 ),
    .din378_WIDTH( 8 ),
    .din379_WIDTH( 8 ),
    .din380_WIDTH( 8 ),
    .din381_WIDTH( 8 ),
    .din382_WIDTH( 8 ),
    .din383_WIDTH( 8 ),
    .din384_WIDTH( 8 ),
    .din385_WIDTH( 8 ),
    .din386_WIDTH( 8 ),
    .din387_WIDTH( 8 ),
    .din388_WIDTH( 8 ),
    .din389_WIDTH( 8 ),
    .din390_WIDTH( 8 ),
    .din391_WIDTH( 8 ),
    .din392_WIDTH( 8 ),
    .din393_WIDTH( 8 ),
    .din394_WIDTH( 8 ),
    .din395_WIDTH( 8 ),
    .din396_WIDTH( 8 ),
    .din397_WIDTH( 8 ),
    .din398_WIDTH( 8 ),
    .din399_WIDTH( 8 ),
    .din400_WIDTH( 8 ),
    .din401_WIDTH( 8 ),
    .din402_WIDTH( 8 ),
    .din403_WIDTH( 8 ),
    .din404_WIDTH( 8 ),
    .din405_WIDTH( 8 ),
    .din406_WIDTH( 8 ),
    .din407_WIDTH( 8 ),
    .din408_WIDTH( 8 ),
    .din409_WIDTH( 8 ),
    .din410_WIDTH( 8 ),
    .din411_WIDTH( 8 ),
    .din412_WIDTH( 8 ),
    .din413_WIDTH( 8 ),
    .din414_WIDTH( 8 ),
    .din415_WIDTH( 8 ),
    .din416_WIDTH( 8 ),
    .din417_WIDTH( 8 ),
    .din418_WIDTH( 8 ),
    .din419_WIDTH( 8 ),
    .din420_WIDTH( 8 ),
    .din421_WIDTH( 8 ),
    .din422_WIDTH( 8 ),
    .din423_WIDTH( 8 ),
    .din424_WIDTH( 8 ),
    .din425_WIDTH( 8 ),
    .din426_WIDTH( 8 ),
    .din427_WIDTH( 8 ),
    .din428_WIDTH( 8 ),
    .din429_WIDTH( 8 ),
    .din430_WIDTH( 8 ),
    .din431_WIDTH( 8 ),
    .din432_WIDTH( 8 ),
    .din433_WIDTH( 8 ),
    .din434_WIDTH( 8 ),
    .din435_WIDTH( 8 ),
    .din436_WIDTH( 8 ),
    .din437_WIDTH( 8 ),
    .din438_WIDTH( 8 ),
    .din439_WIDTH( 8 ),
    .din440_WIDTH( 8 ),
    .din441_WIDTH( 8 ),
    .din442_WIDTH( 8 ),
    .din443_WIDTH( 8 ),
    .din444_WIDTH( 8 ),
    .din445_WIDTH( 8 ),
    .din446_WIDTH( 8 ),
    .din447_WIDTH( 8 ),
    .din448_WIDTH( 8 ),
    .din449_WIDTH( 8 ),
    .din450_WIDTH( 8 ),
    .din451_WIDTH( 8 ),
    .din452_WIDTH( 8 ),
    .din453_WIDTH( 8 ),
    .din454_WIDTH( 8 ),
    .din455_WIDTH( 8 ),
    .din456_WIDTH( 8 ),
    .din457_WIDTH( 8 ),
    .din458_WIDTH( 8 ),
    .din459_WIDTH( 8 ),
    .din460_WIDTH( 8 ),
    .din461_WIDTH( 8 ),
    .din462_WIDTH( 8 ),
    .din463_WIDTH( 8 ),
    .din464_WIDTH( 8 ),
    .din465_WIDTH( 8 ),
    .din466_WIDTH( 8 ),
    .din467_WIDTH( 8 ),
    .din468_WIDTH( 8 ),
    .din469_WIDTH( 8 ),
    .din470_WIDTH( 8 ),
    .din471_WIDTH( 8 ),
    .din472_WIDTH( 8 ),
    .din473_WIDTH( 8 ),
    .din474_WIDTH( 8 ),
    .din475_WIDTH( 8 ),
    .din476_WIDTH( 8 ),
    .din477_WIDTH( 8 ),
    .din478_WIDTH( 8 ),
    .din479_WIDTH( 8 ),
    .din480_WIDTH( 8 ),
    .din481_WIDTH( 8 ),
    .din482_WIDTH( 8 ),
    .din483_WIDTH( 8 ),
    .din484_WIDTH( 8 ),
    .din485_WIDTH( 8 ),
    .din486_WIDTH( 8 ),
    .din487_WIDTH( 8 ),
    .din488_WIDTH( 8 ),
    .din489_WIDTH( 8 ),
    .din490_WIDTH( 8 ),
    .din491_WIDTH( 8 ),
    .din492_WIDTH( 8 ),
    .din493_WIDTH( 8 ),
    .din494_WIDTH( 8 ),
    .din495_WIDTH( 8 ),
    .din496_WIDTH( 8 ),
    .din497_WIDTH( 8 ),
    .din498_WIDTH( 8 ),
    .din499_WIDTH( 8 ),
    .din500_WIDTH( 8 ),
    .din501_WIDTH( 8 ),
    .din502_WIDTH( 8 ),
    .din503_WIDTH( 8 ),
    .din504_WIDTH( 8 ),
    .din505_WIDTH( 8 ),
    .din506_WIDTH( 8 ),
    .din507_WIDTH( 8 ),
    .din508_WIDTH( 8 ),
    .din509_WIDTH( 8 ),
    .din510_WIDTH( 8 ),
    .din511_WIDTH( 8 ),
    .din512_WIDTH( 8 ),
    .din513_WIDTH( 8 ),
    .din514_WIDTH( 8 ),
    .din515_WIDTH( 8 ),
    .din516_WIDTH( 8 ),
    .din517_WIDTH( 8 ),
    .din518_WIDTH( 8 ),
    .din519_WIDTH( 8 ),
    .din520_WIDTH( 8 ),
    .din521_WIDTH( 8 ),
    .din522_WIDTH( 8 ),
    .din523_WIDTH( 8 ),
    .din524_WIDTH( 8 ),
    .din525_WIDTH( 8 ),
    .din526_WIDTH( 8 ),
    .din527_WIDTH( 8 ),
    .din528_WIDTH( 8 ),
    .din529_WIDTH( 8 ),
    .din530_WIDTH( 8 ),
    .din531_WIDTH( 8 ),
    .din532_WIDTH( 8 ),
    .din533_WIDTH( 8 ),
    .din534_WIDTH( 8 ),
    .din535_WIDTH( 8 ),
    .din536_WIDTH( 8 ),
    .din537_WIDTH( 8 ),
    .din538_WIDTH( 8 ),
    .din539_WIDTH( 8 ),
    .din540_WIDTH( 8 ),
    .din541_WIDTH( 8 ),
    .din542_WIDTH( 8 ),
    .din543_WIDTH( 8 ),
    .din544_WIDTH( 8 ),
    .din545_WIDTH( 8 ),
    .din546_WIDTH( 8 ),
    .din547_WIDTH( 8 ),
    .din548_WIDTH( 8 ),
    .din549_WIDTH( 8 ),
    .din550_WIDTH( 8 ),
    .din551_WIDTH( 8 ),
    .din552_WIDTH( 8 ),
    .din553_WIDTH( 8 ),
    .din554_WIDTH( 8 ),
    .din555_WIDTH( 8 ),
    .din556_WIDTH( 8 ),
    .din557_WIDTH( 8 ),
    .din558_WIDTH( 8 ),
    .din559_WIDTH( 8 ),
    .din560_WIDTH( 8 ),
    .din561_WIDTH( 8 ),
    .din562_WIDTH( 8 ),
    .din563_WIDTH( 8 ),
    .din564_WIDTH( 8 ),
    .din565_WIDTH( 8 ),
    .din566_WIDTH( 8 ),
    .din567_WIDTH( 8 ),
    .din568_WIDTH( 8 ),
    .din569_WIDTH( 8 ),
    .din570_WIDTH( 8 ),
    .din571_WIDTH( 8 ),
    .din572_WIDTH( 8 ),
    .din573_WIDTH( 8 ),
    .din574_WIDTH( 8 ),
    .din575_WIDTH( 8 ),
    .din576_WIDTH( 10 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_bkb_U1(
    .din0(tmp_V_fu_1262),
    .din1(tmp_V_1_fu_1266),
    .din2(tmp_V_2_fu_1270),
    .din3(tmp_V_4_fu_1274),
    .din4(tmp_V_5_fu_1278),
    .din5(tmp_V_6_fu_1282),
    .din6(tmp_V_7_fu_1286),
    .din7(tmp_V_8_fu_1290),
    .din8(tmp_V_9_fu_1294),
    .din9(tmp_V_10_fu_1298),
    .din10(tmp_V_11_fu_1302),
    .din11(tmp_V_12_fu_1306),
    .din12(tmp_V_13_fu_1310),
    .din13(tmp_V_14_fu_1314),
    .din14(tmp_V_15_fu_1318),
    .din15(tmp_V_16_fu_1322),
    .din16(tmp_V_17_fu_1326),
    .din17(tmp_V_18_fu_1330),
    .din18(tmp_V_19_fu_1334),
    .din19(tmp_V_20_fu_1338),
    .din20(tmp_V_21_fu_1342),
    .din21(tmp_V_22_fu_1346),
    .din22(tmp_V_23_fu_1350),
    .din23(tmp_V_24_fu_1354),
    .din24(tmp_V_25_fu_1358),
    .din25(tmp_V_26_fu_1362),
    .din26(tmp_V_27_fu_1366),
    .din27(tmp_V_28_fu_1370),
    .din28(tmp_V_29_fu_1374),
    .din29(tmp_V_30_fu_1378),
    .din30(tmp_V_31_fu_1382),
    .din31(tmp_V_32_fu_1386),
    .din32(tmp_V_33_fu_1390),
    .din33(tmp_V_34_fu_1394),
    .din34(tmp_V_35_fu_1398),
    .din35(tmp_V_36_fu_1402),
    .din36(tmp_V_37_fu_1406),
    .din37(tmp_V_38_fu_1410),
    .din38(tmp_V_39_fu_1414),
    .din39(tmp_V_40_fu_1418),
    .din40(tmp_V_41_fu_1422),
    .din41(tmp_V_42_fu_1426),
    .din42(tmp_V_43_fu_1430),
    .din43(tmp_V_44_fu_1434),
    .din44(tmp_V_45_fu_1438),
    .din45(tmp_V_46_fu_1442),
    .din46(tmp_V_47_fu_1446),
    .din47(tmp_V_48_fu_1450),
    .din48(tmp_V_49_fu_1454),
    .din49(tmp_V_50_fu_1458),
    .din50(tmp_V_51_fu_1462),
    .din51(tmp_V_52_fu_1466),
    .din52(tmp_V_53_fu_1470),
    .din53(tmp_V_54_fu_1474),
    .din54(tmp_V_55_fu_1478),
    .din55(tmp_V_56_fu_1482),
    .din56(tmp_V_57_fu_1486),
    .din57(tmp_V_58_fu_1490),
    .din58(tmp_V_59_fu_1494),
    .din59(tmp_V_60_fu_1498),
    .din60(tmp_V_61_fu_1502),
    .din61(tmp_V_62_fu_1506),
    .din62(tmp_V_63_fu_1510),
    .din63(tmp_V_64_fu_1514),
    .din64(tmp_V_65_fu_1518),
    .din65(tmp_V_66_fu_1522),
    .din66(tmp_V_67_fu_1526),
    .din67(tmp_V_68_fu_1530),
    .din68(tmp_V_69_fu_1534),
    .din69(tmp_V_70_fu_1538),
    .din70(tmp_V_71_fu_1542),
    .din71(tmp_V_72_fu_1546),
    .din72(tmp_V_73_fu_1550),
    .din73(tmp_V_74_fu_1554),
    .din74(tmp_V_75_fu_1558),
    .din75(tmp_V_76_fu_1562),
    .din76(tmp_V_77_fu_1566),
    .din77(tmp_V_78_fu_1570),
    .din78(tmp_V_79_fu_1574),
    .din79(tmp_V_80_fu_1578),
    .din80(tmp_V_81_fu_1582),
    .din81(tmp_V_82_fu_1586),
    .din82(tmp_V_83_fu_1590),
    .din83(tmp_V_84_fu_1594),
    .din84(tmp_V_85_fu_1598),
    .din85(tmp_V_86_fu_1602),
    .din86(tmp_V_87_fu_1606),
    .din87(tmp_V_88_fu_1610),
    .din88(tmp_V_89_fu_1614),
    .din89(tmp_V_90_fu_1618),
    .din90(tmp_V_91_fu_1622),
    .din91(tmp_V_92_fu_1626),
    .din92(tmp_V_93_fu_1630),
    .din93(tmp_V_94_fu_1634),
    .din94(tmp_V_95_fu_1638),
    .din95(tmp_V_96_fu_1642),
    .din96(tmp_V_97_fu_1646),
    .din97(tmp_V_98_fu_1650),
    .din98(tmp_V_99_fu_1654),
    .din99(tmp_V_100_fu_1658),
    .din100(tmp_V_101_fu_1662),
    .din101(tmp_V_102_fu_1666),
    .din102(tmp_V_103_fu_1670),
    .din103(tmp_V_104_fu_1674),
    .din104(tmp_V_105_fu_1678),
    .din105(tmp_V_106_fu_1682),
    .din106(tmp_V_107_fu_1686),
    .din107(tmp_V_108_fu_1690),
    .din108(tmp_V_109_fu_1694),
    .din109(tmp_V_110_fu_1698),
    .din110(tmp_V_111_fu_1702),
    .din111(tmp_V_112_fu_1706),
    .din112(tmp_V_113_fu_1710),
    .din113(tmp_V_114_fu_1714),
    .din114(tmp_V_115_fu_1718),
    .din115(tmp_V_116_fu_1722),
    .din116(tmp_V_117_fu_1726),
    .din117(tmp_V_118_fu_1730),
    .din118(tmp_V_119_fu_1734),
    .din119(tmp_V_120_fu_1738),
    .din120(tmp_V_121_fu_1742),
    .din121(tmp_V_122_fu_1746),
    .din122(tmp_V_123_fu_1750),
    .din123(tmp_V_124_fu_1754),
    .din124(tmp_V_125_fu_1758),
    .din125(tmp_V_126_fu_1762),
    .din126(tmp_V_127_fu_1766),
    .din127(tmp_V_128_fu_1770),
    .din128(tmp_V_129_fu_1774),
    .din129(tmp_V_130_fu_1778),
    .din130(tmp_V_131_fu_1782),
    .din131(tmp_V_132_fu_1786),
    .din132(tmp_V_133_fu_1790),
    .din133(tmp_V_134_fu_1794),
    .din134(tmp_V_135_fu_1798),
    .din135(tmp_V_136_fu_1802),
    .din136(tmp_V_137_fu_1806),
    .din137(tmp_V_138_fu_1810),
    .din138(tmp_V_139_fu_1814),
    .din139(tmp_V_140_fu_1818),
    .din140(tmp_V_141_fu_1822),
    .din141(tmp_V_142_fu_1826),
    .din142(tmp_V_143_fu_1830),
    .din143(tmp_V_144_fu_1834),
    .din144(tmp_V_145_fu_1838),
    .din145(tmp_V_146_fu_1842),
    .din146(tmp_V_147_fu_1846),
    .din147(tmp_V_148_fu_1850),
    .din148(tmp_V_149_fu_1854),
    .din149(tmp_V_150_fu_1858),
    .din150(tmp_V_151_fu_1862),
    .din151(tmp_V_152_fu_1866),
    .din152(tmp_V_153_fu_1870),
    .din153(tmp_V_154_fu_1874),
    .din154(tmp_V_155_fu_1878),
    .din155(tmp_V_156_fu_1882),
    .din156(tmp_V_157_fu_1886),
    .din157(tmp_V_158_fu_1890),
    .din158(tmp_V_159_fu_1894),
    .din159(tmp_V_160_fu_1898),
    .din160(tmp_V_161_fu_1902),
    .din161(tmp_V_162_fu_1906),
    .din162(tmp_V_163_fu_1910),
    .din163(tmp_V_164_fu_1914),
    .din164(tmp_V_165_fu_1918),
    .din165(tmp_V_166_fu_1922),
    .din166(tmp_V_167_fu_1926),
    .din167(tmp_V_168_fu_1930),
    .din168(tmp_V_169_fu_1934),
    .din169(tmp_V_170_fu_1938),
    .din170(tmp_V_171_fu_1942),
    .din171(tmp_V_172_fu_1946),
    .din172(tmp_V_173_fu_1950),
    .din173(tmp_V_174_fu_1954),
    .din174(tmp_V_175_fu_1958),
    .din175(tmp_V_176_fu_1962),
    .din176(tmp_V_177_fu_1966),
    .din177(tmp_V_178_fu_1970),
    .din178(tmp_V_179_fu_1974),
    .din179(tmp_V_180_fu_1978),
    .din180(tmp_V_181_fu_1982),
    .din181(tmp_V_182_fu_1986),
    .din182(tmp_V_183_fu_1990),
    .din183(tmp_V_184_fu_1994),
    .din184(tmp_V_185_fu_1998),
    .din185(tmp_V_186_fu_2002),
    .din186(tmp_V_187_fu_2006),
    .din187(tmp_V_188_fu_2010),
    .din188(tmp_V_189_fu_2014),
    .din189(tmp_V_190_fu_2018),
    .din190(tmp_V_191_fu_2022),
    .din191(tmp_V_192_fu_2026),
    .din192(tmp_V_193_fu_2030),
    .din193(tmp_V_194_fu_2034),
    .din194(tmp_V_195_fu_2038),
    .din195(tmp_V_196_fu_2042),
    .din196(tmp_V_197_fu_2046),
    .din197(tmp_V_198_fu_2050),
    .din198(tmp_V_199_fu_2054),
    .din199(tmp_V_200_fu_2058),
    .din200(tmp_V_201_fu_2062),
    .din201(tmp_V_202_fu_2066),
    .din202(tmp_V_203_fu_2070),
    .din203(tmp_V_204_fu_2074),
    .din204(tmp_V_205_fu_2078),
    .din205(tmp_V_206_fu_2082),
    .din206(tmp_V_207_fu_2086),
    .din207(tmp_V_208_fu_2090),
    .din208(tmp_V_209_fu_2094),
    .din209(tmp_V_210_fu_2098),
    .din210(tmp_V_211_fu_2102),
    .din211(tmp_V_212_fu_2106),
    .din212(tmp_V_213_fu_2110),
    .din213(tmp_V_214_fu_2114),
    .din214(tmp_V_215_fu_2118),
    .din215(tmp_V_216_fu_2122),
    .din216(tmp_V_217_fu_2126),
    .din217(tmp_V_218_fu_2130),
    .din218(tmp_V_219_fu_2134),
    .din219(tmp_V_220_fu_2138),
    .din220(tmp_V_221_fu_2142),
    .din221(tmp_V_222_fu_2146),
    .din222(tmp_V_223_fu_2150),
    .din223(tmp_V_224_fu_2154),
    .din224(tmp_V_225_fu_2158),
    .din225(tmp_V_226_fu_2162),
    .din226(tmp_V_227_fu_2166),
    .din227(tmp_V_228_fu_2170),
    .din228(tmp_V_229_fu_2174),
    .din229(tmp_V_230_fu_2178),
    .din230(tmp_V_231_fu_2182),
    .din231(tmp_V_232_fu_2186),
    .din232(tmp_V_233_fu_2190),
    .din233(tmp_V_234_fu_2194),
    .din234(tmp_V_235_fu_2198),
    .din235(tmp_V_236_fu_2202),
    .din236(tmp_V_237_fu_2206),
    .din237(tmp_V_238_fu_2210),
    .din238(tmp_V_239_fu_2214),
    .din239(tmp_V_240_fu_2218),
    .din240(tmp_V_241_fu_2222),
    .din241(tmp_V_242_fu_2226),
    .din242(tmp_V_243_fu_2230),
    .din243(tmp_V_244_fu_2234),
    .din244(tmp_V_245_fu_2238),
    .din245(tmp_V_246_fu_2242),
    .din246(tmp_V_247_fu_2246),
    .din247(tmp_V_248_fu_2250),
    .din248(tmp_V_249_fu_2254),
    .din249(tmp_V_250_fu_2258),
    .din250(tmp_V_251_fu_2262),
    .din251(tmp_V_252_fu_2266),
    .din252(tmp_V_253_fu_2270),
    .din253(tmp_V_254_fu_2274),
    .din254(tmp_V_255_fu_2278),
    .din255(tmp_V_256_fu_2282),
    .din256(tmp_V_257_fu_2286),
    .din257(tmp_V_258_fu_2290),
    .din258(tmp_V_259_fu_2294),
    .din259(tmp_V_260_fu_2298),
    .din260(tmp_V_261_fu_2302),
    .din261(tmp_V_262_fu_2306),
    .din262(tmp_V_263_fu_2310),
    .din263(tmp_V_264_fu_2314),
    .din264(tmp_V_265_fu_2318),
    .din265(tmp_V_266_fu_2322),
    .din266(tmp_V_267_fu_2326),
    .din267(tmp_V_268_fu_2330),
    .din268(tmp_V_269_fu_2334),
    .din269(tmp_V_270_fu_2338),
    .din270(tmp_V_271_fu_2342),
    .din271(tmp_V_272_fu_2346),
    .din272(tmp_V_273_fu_2350),
    .din273(tmp_V_274_fu_2354),
    .din274(tmp_V_275_fu_2358),
    .din275(tmp_V_276_fu_2362),
    .din276(tmp_V_277_fu_2366),
    .din277(tmp_V_278_fu_2370),
    .din278(tmp_V_279_fu_2374),
    .din279(tmp_V_280_fu_2378),
    .din280(tmp_V_281_fu_2382),
    .din281(tmp_V_282_fu_2386),
    .din282(tmp_V_283_fu_2390),
    .din283(tmp_V_284_fu_2394),
    .din284(tmp_V_285_fu_2398),
    .din285(tmp_V_286_fu_2402),
    .din286(tmp_V_287_fu_2406),
    .din287(tmp_V_288_fu_2410),
    .din288(tmp_V_289_fu_2414),
    .din289(tmp_V_290_fu_2418),
    .din290(tmp_V_291_fu_2422),
    .din291(tmp_V_292_fu_2426),
    .din292(tmp_V_293_fu_2430),
    .din293(tmp_V_294_fu_2434),
    .din294(tmp_V_295_fu_2438),
    .din295(tmp_V_296_fu_2442),
    .din296(tmp_V_297_fu_2446),
    .din297(tmp_V_298_fu_2450),
    .din298(tmp_V_299_fu_2454),
    .din299(tmp_V_300_fu_2458),
    .din300(tmp_V_301_fu_2462),
    .din301(tmp_V_302_fu_2466),
    .din302(tmp_V_303_fu_2470),
    .din303(tmp_V_304_fu_2474),
    .din304(tmp_V_305_fu_2478),
    .din305(tmp_V_306_fu_2482),
    .din306(tmp_V_307_fu_2486),
    .din307(tmp_V_308_fu_2490),
    .din308(tmp_V_309_fu_2494),
    .din309(tmp_V_310_fu_2498),
    .din310(tmp_V_311_fu_2502),
    .din311(tmp_V_312_fu_2506),
    .din312(tmp_V_313_fu_2510),
    .din313(tmp_V_314_fu_2514),
    .din314(tmp_V_315_fu_2518),
    .din315(tmp_V_316_fu_2522),
    .din316(tmp_V_317_fu_2526),
    .din317(tmp_V_318_fu_2530),
    .din318(tmp_V_319_fu_2534),
    .din319(tmp_V_320_fu_2538),
    .din320(tmp_V_321_fu_2542),
    .din321(tmp_V_322_fu_2546),
    .din322(tmp_V_323_fu_2550),
    .din323(tmp_V_324_fu_2554),
    .din324(tmp_V_325_fu_2558),
    .din325(tmp_V_326_fu_2562),
    .din326(tmp_V_327_fu_2566),
    .din327(tmp_V_328_fu_2570),
    .din328(tmp_V_329_fu_2574),
    .din329(tmp_V_330_fu_2578),
    .din330(tmp_V_331_fu_2582),
    .din331(tmp_V_332_fu_2586),
    .din332(tmp_V_333_fu_2590),
    .din333(tmp_V_334_fu_2594),
    .din334(tmp_V_335_fu_2598),
    .din335(tmp_V_336_fu_2602),
    .din336(tmp_V_337_fu_2606),
    .din337(tmp_V_338_fu_2610),
    .din338(tmp_V_339_fu_2614),
    .din339(tmp_V_340_fu_2618),
    .din340(tmp_V_341_fu_2622),
    .din341(tmp_V_342_fu_2626),
    .din342(tmp_V_343_fu_2630),
    .din343(tmp_V_344_fu_2634),
    .din344(tmp_V_345_fu_2638),
    .din345(tmp_V_346_fu_2642),
    .din346(tmp_V_347_fu_2646),
    .din347(tmp_V_348_fu_2650),
    .din348(tmp_V_349_fu_2654),
    .din349(tmp_V_350_fu_2658),
    .din350(tmp_V_351_fu_2662),
    .din351(tmp_V_352_fu_2666),
    .din352(tmp_V_353_fu_2670),
    .din353(tmp_V_354_fu_2674),
    .din354(tmp_V_355_fu_2678),
    .din355(tmp_V_356_fu_2682),
    .din356(tmp_V_357_fu_2686),
    .din357(tmp_V_358_fu_2690),
    .din358(tmp_V_359_fu_2694),
    .din359(tmp_V_360_fu_2698),
    .din360(tmp_V_361_fu_2702),
    .din361(tmp_V_362_fu_2706),
    .din362(tmp_V_363_fu_2710),
    .din363(tmp_V_364_fu_2714),
    .din364(tmp_V_365_fu_2718),
    .din365(tmp_V_366_fu_2722),
    .din366(tmp_V_367_fu_2726),
    .din367(tmp_V_368_fu_2730),
    .din368(tmp_V_369_fu_2734),
    .din369(tmp_V_370_fu_2738),
    .din370(tmp_V_371_fu_2742),
    .din371(tmp_V_372_fu_2746),
    .din372(tmp_V_373_fu_2750),
    .din373(tmp_V_374_fu_2754),
    .din374(tmp_V_375_fu_2758),
    .din375(tmp_V_376_fu_2762),
    .din376(tmp_V_377_fu_2766),
    .din377(tmp_V_378_fu_2770),
    .din378(tmp_V_379_fu_2774),
    .din379(tmp_V_380_fu_2778),
    .din380(tmp_V_381_fu_2782),
    .din381(tmp_V_382_fu_2786),
    .din382(tmp_V_383_fu_2790),
    .din383(tmp_V_384_fu_2794),
    .din384(tmp_V_385_fu_2798),
    .din385(tmp_V_386_fu_2802),
    .din386(tmp_V_387_fu_2806),
    .din387(tmp_V_388_fu_2810),
    .din388(tmp_V_389_fu_2814),
    .din389(tmp_V_390_fu_2818),
    .din390(tmp_V_391_fu_2822),
    .din391(tmp_V_392_fu_2826),
    .din392(tmp_V_393_fu_2830),
    .din393(tmp_V_394_fu_2834),
    .din394(tmp_V_395_fu_2838),
    .din395(tmp_V_396_fu_2842),
    .din396(tmp_V_397_fu_2846),
    .din397(tmp_V_398_fu_2850),
    .din398(tmp_V_399_fu_2854),
    .din399(tmp_V_400_fu_2858),
    .din400(tmp_V_401_fu_2862),
    .din401(tmp_V_402_fu_2866),
    .din402(tmp_V_403_fu_2870),
    .din403(tmp_V_404_fu_2874),
    .din404(tmp_V_405_fu_2878),
    .din405(tmp_V_406_fu_2882),
    .din406(tmp_V_407_fu_2886),
    .din407(tmp_V_408_fu_2890),
    .din408(tmp_V_409_fu_2894),
    .din409(tmp_V_410_fu_2898),
    .din410(tmp_V_411_fu_2902),
    .din411(tmp_V_412_fu_2906),
    .din412(tmp_V_413_fu_2910),
    .din413(tmp_V_414_fu_2914),
    .din414(tmp_V_415_fu_2918),
    .din415(tmp_V_416_fu_2922),
    .din416(tmp_V_417_fu_2926),
    .din417(tmp_V_418_fu_2930),
    .din418(tmp_V_419_fu_2934),
    .din419(tmp_V_420_fu_2938),
    .din420(tmp_V_421_fu_2942),
    .din421(tmp_V_422_fu_2946),
    .din422(tmp_V_423_fu_2950),
    .din423(tmp_V_424_fu_2954),
    .din424(tmp_V_425_fu_2958),
    .din425(tmp_V_426_fu_2962),
    .din426(tmp_V_427_fu_2966),
    .din427(tmp_V_428_fu_2970),
    .din428(tmp_V_429_fu_2974),
    .din429(tmp_V_430_fu_2978),
    .din430(tmp_V_431_fu_2982),
    .din431(tmp_V_432_fu_2986),
    .din432(tmp_V_433_fu_2990),
    .din433(tmp_V_434_fu_2994),
    .din434(tmp_V_435_fu_2998),
    .din435(tmp_V_436_fu_3002),
    .din436(tmp_V_437_fu_3006),
    .din437(tmp_V_438_fu_3010),
    .din438(tmp_V_439_fu_3014),
    .din439(tmp_V_440_fu_3018),
    .din440(tmp_V_441_fu_3022),
    .din441(tmp_V_442_fu_3026),
    .din442(tmp_V_443_fu_3030),
    .din443(tmp_V_444_fu_3034),
    .din444(tmp_V_445_fu_3038),
    .din445(tmp_V_446_fu_3042),
    .din446(tmp_V_447_fu_3046),
    .din447(tmp_V_448_fu_3050),
    .din448(tmp_V_449_fu_3054),
    .din449(tmp_V_450_fu_3058),
    .din450(tmp_V_451_fu_3062),
    .din451(tmp_V_452_fu_3066),
    .din452(tmp_V_453_fu_3070),
    .din453(tmp_V_454_fu_3074),
    .din454(tmp_V_455_fu_3078),
    .din455(tmp_V_456_fu_3082),
    .din456(tmp_V_457_fu_3086),
    .din457(tmp_V_458_fu_3090),
    .din458(tmp_V_459_fu_3094),
    .din459(tmp_V_460_fu_3098),
    .din460(tmp_V_461_fu_3102),
    .din461(tmp_V_462_fu_3106),
    .din462(tmp_V_463_fu_3110),
    .din463(tmp_V_464_fu_3114),
    .din464(tmp_V_465_fu_3118),
    .din465(tmp_V_466_fu_3122),
    .din466(tmp_V_467_fu_3126),
    .din467(tmp_V_468_fu_3130),
    .din468(tmp_V_469_fu_3134),
    .din469(tmp_V_470_fu_3138),
    .din470(tmp_V_471_fu_3142),
    .din471(tmp_V_472_fu_3146),
    .din472(tmp_V_473_fu_3150),
    .din473(tmp_V_474_fu_3154),
    .din474(tmp_V_475_fu_3158),
    .din475(tmp_V_476_fu_3162),
    .din476(tmp_V_477_fu_3166),
    .din477(tmp_V_478_fu_3170),
    .din478(tmp_V_479_fu_3174),
    .din479(tmp_V_480_fu_3178),
    .din480(tmp_V_481_fu_3182),
    .din481(tmp_V_482_fu_3186),
    .din482(tmp_V_483_fu_3190),
    .din483(tmp_V_484_fu_3194),
    .din484(tmp_V_485_fu_3198),
    .din485(tmp_V_486_fu_3202),
    .din486(tmp_V_487_fu_3206),
    .din487(tmp_V_488_fu_3210),
    .din488(tmp_V_489_fu_3214),
    .din489(tmp_V_490_fu_3218),
    .din490(tmp_V_491_fu_3222),
    .din491(tmp_V_492_fu_3226),
    .din492(tmp_V_493_fu_3230),
    .din493(tmp_V_494_fu_3234),
    .din494(tmp_V_495_fu_3238),
    .din495(tmp_V_496_fu_3242),
    .din496(tmp_V_497_fu_3246),
    .din497(tmp_V_498_fu_3250),
    .din498(tmp_V_499_fu_3254),
    .din499(tmp_V_500_fu_3258),
    .din500(tmp_V_501_fu_3262),
    .din501(tmp_V_502_fu_3266),
    .din502(tmp_V_503_fu_3270),
    .din503(tmp_V_504_fu_3274),
    .din504(tmp_V_505_fu_3278),
    .din505(tmp_V_506_fu_3282),
    .din506(tmp_V_507_fu_3286),
    .din507(tmp_V_508_fu_3290),
    .din508(tmp_V_509_fu_3294),
    .din509(tmp_V_510_fu_3298),
    .din510(tmp_V_511_fu_3302),
    .din511(tmp_V_512_fu_3306),
    .din512(tmp_V_513_fu_3310),
    .din513(tmp_V_514_fu_3314),
    .din514(tmp_V_515_fu_3318),
    .din515(tmp_V_516_fu_3322),
    .din516(tmp_V_517_fu_3326),
    .din517(tmp_V_518_fu_3330),
    .din518(tmp_V_519_fu_3334),
    .din519(tmp_V_520_fu_3338),
    .din520(tmp_V_521_fu_3342),
    .din521(tmp_V_522_fu_3346),
    .din522(tmp_V_523_fu_3350),
    .din523(tmp_V_524_fu_3354),
    .din524(tmp_V_525_fu_3358),
    .din525(tmp_V_526_fu_3362),
    .din526(tmp_V_527_fu_3366),
    .din527(tmp_V_528_fu_3370),
    .din528(tmp_V_529_fu_3374),
    .din529(tmp_V_530_fu_3378),
    .din530(tmp_V_531_fu_3382),
    .din531(tmp_V_532_fu_3386),
    .din532(tmp_V_533_fu_3390),
    .din533(tmp_V_534_fu_3394),
    .din534(tmp_V_535_fu_3398),
    .din535(tmp_V_536_fu_3402),
    .din536(tmp_V_537_fu_3406),
    .din537(tmp_V_538_fu_3410),
    .din538(tmp_V_539_fu_3414),
    .din539(tmp_V_540_fu_3418),
    .din540(tmp_V_541_fu_3422),
    .din541(tmp_V_542_fu_3426),
    .din542(tmp_V_543_fu_3430),
    .din543(tmp_V_544_fu_3434),
    .din544(tmp_V_545_fu_3438),
    .din545(tmp_V_546_fu_3442),
    .din546(tmp_V_547_fu_3446),
    .din547(tmp_V_548_fu_3450),
    .din548(tmp_V_549_fu_3454),
    .din549(tmp_V_550_fu_3458),
    .din550(tmp_V_551_fu_3462),
    .din551(tmp_V_552_fu_3466),
    .din552(tmp_V_553_fu_3470),
    .din553(tmp_V_554_fu_3474),
    .din554(tmp_V_555_fu_3478),
    .din555(tmp_V_556_fu_3482),
    .din556(tmp_V_557_fu_3486),
    .din557(tmp_V_558_fu_3490),
    .din558(tmp_V_559_fu_3494),
    .din559(tmp_V_560_fu_3498),
    .din560(tmp_V_561_fu_3502),
    .din561(tmp_V_562_fu_3506),
    .din562(tmp_V_563_fu_3510),
    .din563(tmp_V_564_fu_3514),
    .din564(tmp_V_565_fu_3518),
    .din565(tmp_V_566_fu_3522),
    .din566(tmp_V_567_fu_3526),
    .din567(tmp_V_568_fu_3530),
    .din568(tmp_V_569_fu_3534),
    .din569(tmp_V_570_fu_3538),
    .din570(tmp_V_571_fu_3542),
    .din571(tmp_V_572_fu_3546),
    .din572(tmp_V_573_fu_3550),
    .din573(tmp_V_574_fu_3554),
    .din574(tmp_V_575_fu_3558),
    .din575(tmp_V_576_fu_3562),
    .din576(inElem_V_1_fu_6525_p577),
    .dout(inElem_V_1_fu_6525_p578)
);

StreamingFCLayer_Batch_0_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U2(
    .din0(mul_ln1352_fu_10718_p0),
    .din1(trunc_ln647_reg_15064),
    .dout(mul_ln1352_fu_10718_p2)
);

StreamingFCLayer_Batch_0_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U3(
    .din0(mul_ln1352_1_fu_10745_p0),
    .din1(p_Result_1_0_1_reg_15069),
    .dout(mul_ln1352_1_fu_10745_p2)
);

StreamingFCLayer_Batch_0_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U4(
    .din0(mul_ln1352_2_fu_10774_p0),
    .din1(p_Result_1_1_reg_15074),
    .dout(mul_ln1352_2_fu_10774_p2)
);

StreamingFCLayer_Batch_0_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U5(
    .din0(mul_ln1352_3_fu_10787_p0),
    .din1(p_Result_1_1_1_reg_15079),
    .dout(mul_ln1352_3_fu_10787_p2)
);

StreamingFCLayer_Batch_0_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U6(
    .din0(mul_ln1352_4_fu_10816_p0),
    .din1(p_Result_1_2_reg_15084),
    .dout(mul_ln1352_4_fu_10816_p2)
);

StreamingFCLayer_Batch_0_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U7(
    .din0(mul_ln1352_5_fu_10829_p0),
    .din1(p_Result_1_2_1_reg_15089),
    .dout(mul_ln1352_5_fu_10829_p2)
);

StreamingFCLayer_Batch_0_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U8(
    .din0(mul_ln1352_6_fu_10858_p0),
    .din1(p_Result_1_3_reg_15094),
    .dout(mul_ln1352_6_fu_10858_p2)
);

StreamingFCLayer_Batch_0_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U9(
    .din0(mul_ln1352_7_fu_10871_p0),
    .din1(p_Result_1_3_1_reg_15099),
    .dout(mul_ln1352_7_fu_10871_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd0) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_3600 <= inElem_V_1_fu_6525_p578;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd214)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd213)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd212)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd211)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd210)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd209)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd208)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd207)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd206)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd205)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd204)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd203)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd202)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd201)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd200)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd199)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd198)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd197)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd196)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd195)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd194)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd193)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd192)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd191)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd190)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd189)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd188)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd187)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd186)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd185)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd184)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd183)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd182)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd181)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd180)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd179)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd178)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd177)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd176)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd175)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd174)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd173)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd172)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd171)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd170)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd169)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd168)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd167)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd166)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd165)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd164)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd163)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd162)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd161)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd160)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd159)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd158)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd157)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd156)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd155)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd154)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd153)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd152)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd151)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd150)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd149)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd148)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd147)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd146)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd145)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd144)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd143)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd142)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd141)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd140)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd139)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd138)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd137)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd136)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd135)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd134)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd133)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd132)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd131)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd130)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd129)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd128)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd127)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd126)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd125)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd124)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd123)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd122)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd121)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd120)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd119)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd118)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd117)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd116)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd115)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd114)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd113)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd112)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd111)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd110)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd109)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd108)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd107)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd106)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd105)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd104)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd103)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd102)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd101)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd100)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd99)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd98)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd97)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd96)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd95)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd94)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd93)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd92)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd91)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd90)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd89)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd88)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd87)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd86)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd85)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd84)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd83)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd82)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd81)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd80)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd79)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd78)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd77)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd76)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd75)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd74)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd73)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd72)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd71)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd70)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd69)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd68)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd67)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd66)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd65)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd64)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd63)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd62)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd61)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd60)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd59)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd58)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd57)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd56)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd55)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd54)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd53)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd52)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd51)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd50)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd49)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd48)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd47)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd46)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd45)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd44)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd43)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd42)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd41)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd40)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd39)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd38)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd37)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd36)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd35)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd34)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd33)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd32)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd31)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd30)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd29)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd28)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd27)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd26)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd574)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd573)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd572)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd25)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd571)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd570)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd569)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd568)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd567)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd566)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd565)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd564)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd563)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd562)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd24)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd561)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd560)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd559)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd558)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd557)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd556)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd555)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd554)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd553)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd552)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd23)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd551)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd550)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd549)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd548)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd547)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd546)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd545)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd544)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd543)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd542)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd22)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd541)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd540)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd539)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd538)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd537)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd536)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd535)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd534)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd533)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd532)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd21)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd531)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd530)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd529)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd528)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd527)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd526)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd525)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd524)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd523)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd522)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd20)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd521)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd520)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd519)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd518)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd517)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd516)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd515)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd514)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd513)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd512)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd19)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd511)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd510)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd509)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd508)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd507)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd506)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd505)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd504)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd503)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd502)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd18)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd501)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd500)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd499)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd498)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd497)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd496)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd495)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd494)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd493)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd492)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd17)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd491)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd490)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd489)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd488)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd487)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd486)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd485)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd484)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd483)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd482)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd16)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd481)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd480)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd479)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd478)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd477)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd476)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd475)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd474)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd473)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd472)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd15)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd471)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd470)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd469)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd468)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd467)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd466)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd465)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd464)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd463)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd462)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd14)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd461)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd460)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd459)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd458)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd457)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd456)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd455)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd454)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd453)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd452)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd13)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd451)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd450)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd449)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd448)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd447)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd446)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd445)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd444)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd443)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd442)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd12)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd441)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd440)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd439)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd438)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd437)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd436)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd435)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd434)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd433)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd432)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd11)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd431)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd430)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd429)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd428)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd427)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd426)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd425)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd424)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd423)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd422)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd10)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd421)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd420)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd419)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd418)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd417)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd416)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd415)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd414)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd413)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd412)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd9)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd411)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd410)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd409)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd408)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd407)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd406)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd405)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd404)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd403)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd402)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd8)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd401)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd400)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd399)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd398)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd397)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd396)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd395)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd394)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd393)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd392)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd7)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd391)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd390)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd389)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd388)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd387)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd386)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd385)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd384)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd383)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd382)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd6)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd381)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd380)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd379)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd378)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd377)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd376)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd375)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd374)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd373)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd372)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd5)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd371)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd370)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd369)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd368)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd367)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd366)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd365)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd364)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd363)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd362)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd4)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd361)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd360)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd359)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd358)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd357)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd356)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd355)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd354)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd353)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd352)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd3)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd351)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd350)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd349)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd348)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd347)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd346)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd345)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd344)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd343)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd342)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd2)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd341)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd340)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd339)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd338)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd337)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd336)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd335)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd334)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd333)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd332)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd331)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd330)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd329)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd328)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd327)) | (~(trunc_ln321_fu_7683_p1 == 10'd214) & ~(trunc_ln321_fu_7683_p1 == 10'd213) & ~(trunc_ln321_fu_7683_p1 == 10'd212) & ~(trunc_ln321_fu_7683_p1 == 10'd211) & ~(trunc_ln321_fu_7683_p1 == 10'd210) & ~(trunc_ln321_fu_7683_p1 == 10'd209) & ~(trunc_ln321_fu_7683_p1 == 10'd208) & ~(trunc_ln321_fu_7683_p1 == 10'd207) & ~(trunc_ln321_fu_7683_p1 == 10'd206) & ~(trunc_ln321_fu_7683_p1 == 10'd205) & ~(trunc_ln321_fu_7683_p1 == 10'd204) & ~(trunc_ln321_fu_7683_p1 == 10'd203) & ~(trunc_ln321_fu_7683_p1 == 10'd202) & ~(trunc_ln321_fu_7683_p1 == 10'd201) & ~(trunc_ln321_fu_7683_p1 == 10'd200) & ~(trunc_ln321_fu_7683_p1 == 10'd199) & ~(trunc_ln321_fu_7683_p1 == 10'd198) & ~(trunc_ln321_fu_7683_p1 == 10'd197) & ~(trunc_ln321_fu_7683_p1 == 10'd196) & ~(trunc_ln321_fu_7683_p1 == 10'd195) & ~(trunc_ln321_fu_7683_p1 == 10'd194) & ~(trunc_ln321_fu_7683_p1 == 10'd193) & ~(trunc_ln321_fu_7683_p1 == 10'd192) & ~(trunc_ln321_fu_7683_p1 == 10'd191) & ~(trunc_ln321_fu_7683_p1 == 10'd190) & ~(trunc_ln321_fu_7683_p1 == 10'd189) & ~(trunc_ln321_fu_7683_p1 == 10'd188) & ~(trunc_ln321_fu_7683_p1 == 10'd187) & ~(trunc_ln321_fu_7683_p1 == 10'd186) & ~(trunc_ln321_fu_7683_p1 == 10'd185) & ~(trunc_ln321_fu_7683_p1 == 10'd184) & ~(trunc_ln321_fu_7683_p1 == 10'd183) & ~(trunc_ln321_fu_7683_p1 == 10'd182) & ~(trunc_ln321_fu_7683_p1 == 10'd181) & ~(trunc_ln321_fu_7683_p1 == 10'd180) & ~(trunc_ln321_fu_7683_p1 == 10'd179) & ~(trunc_ln321_fu_7683_p1 == 10'd178) & ~(trunc_ln321_fu_7683_p1 == 10'd177) & ~(trunc_ln321_fu_7683_p1 == 10'd176) & ~(trunc_ln321_fu_7683_p1 == 10'd175) & ~(trunc_ln321_fu_7683_p1 == 10'd174) & ~(trunc_ln321_fu_7683_p1 == 10'd173) & ~(trunc_ln321_fu_7683_p1 == 10'd172) & ~(trunc_ln321_fu_7683_p1 == 10'd171) & ~(trunc_ln321_fu_7683_p1 == 10'd170) & ~(trunc_ln321_fu_7683_p1 == 10'd169) & ~(trunc_ln321_fu_7683_p1 == 10'd168) & ~(trunc_ln321_fu_7683_p1 == 10'd167) & ~(trunc_ln321_fu_7683_p1 == 10'd166) & ~(trunc_ln321_fu_7683_p1 == 10'd165) & ~(trunc_ln321_fu_7683_p1 == 10'd164) & ~(trunc_ln321_fu_7683_p1 == 10'd163) & ~(trunc_ln321_fu_7683_p1 == 10'd162) & ~(trunc_ln321_fu_7683_p1 == 10'd161) & ~(trunc_ln321_fu_7683_p1 == 10'd160) & ~(trunc_ln321_fu_7683_p1 == 10'd159) & ~(trunc_ln321_fu_7683_p1 == 10'd158) & ~(trunc_ln321_fu_7683_p1 == 10'd157) & ~(trunc_ln321_fu_7683_p1 == 10'd156) & ~(trunc_ln321_fu_7683_p1 == 10'd155) & ~(trunc_ln321_fu_7683_p1 == 10'd154) & ~(trunc_ln321_fu_7683_p1 == 10'd153) & ~(trunc_ln321_fu_7683_p1 == 10'd152) & ~(trunc_ln321_fu_7683_p1 == 10'd151) & ~(trunc_ln321_fu_7683_p1 == 10'd150) & ~(trunc_ln321_fu_7683_p1 == 10'd149) & ~(trunc_ln321_fu_7683_p1 == 10'd148) & ~(trunc_ln321_fu_7683_p1 == 10'd147) & ~(trunc_ln321_fu_7683_p1 == 10'd146) & ~(trunc_ln321_fu_7683_p1 == 10'd145) & ~(trunc_ln321_fu_7683_p1 == 10'd144) & ~(trunc_ln321_fu_7683_p1 == 10'd143) & ~(trunc_ln321_fu_7683_p1 == 10'd142) & ~(trunc_ln321_fu_7683_p1 == 10'd141) & ~(trunc_ln321_fu_7683_p1 == 10'd140) & ~(trunc_ln321_fu_7683_p1 == 10'd139) & ~(trunc_ln321_fu_7683_p1 == 10'd138) & ~(trunc_ln321_fu_7683_p1 == 10'd137) & ~(trunc_ln321_fu_7683_p1 == 10'd136) & ~(trunc_ln321_fu_7683_p1 == 10'd135) & ~(trunc_ln321_fu_7683_p1 == 10'd134) & ~(trunc_ln321_fu_7683_p1 == 10'd133) & ~(trunc_ln321_fu_7683_p1 == 10'd132) & ~(trunc_ln321_fu_7683_p1 == 10'd131) & ~(trunc_ln321_fu_7683_p1 == 10'd130) & ~(trunc_ln321_fu_7683_p1 == 10'd129) & ~(trunc_ln321_fu_7683_p1 == 10'd128) & ~(trunc_ln321_fu_7683_p1 == 10'd127) & ~(trunc_ln321_fu_7683_p1 == 10'd126) & ~(trunc_ln321_fu_7683_p1 == 10'd125) & ~(trunc_ln321_fu_7683_p1 == 10'd124) & ~(trunc_ln321_fu_7683_p1 == 10'd123) & ~(trunc_ln321_fu_7683_p1 == 10'd122) & ~(trunc_ln321_fu_7683_p1 == 10'd121) & ~(trunc_ln321_fu_7683_p1 == 10'd120) & ~(trunc_ln321_fu_7683_p1 == 10'd119) & ~(trunc_ln321_fu_7683_p1 == 10'd118) & ~(trunc_ln321_fu_7683_p1 == 10'd117) & ~(trunc_ln321_fu_7683_p1 == 10'd116) & ~(trunc_ln321_fu_7683_p1 == 10'd115) & ~(trunc_ln321_fu_7683_p1 == 10'd114) & ~(trunc_ln321_fu_7683_p1 == 10'd113) & ~(trunc_ln321_fu_7683_p1 == 10'd112) & ~(trunc_ln321_fu_7683_p1 == 10'd111) & ~(trunc_ln321_fu_7683_p1 == 10'd110) & ~(trunc_ln321_fu_7683_p1 == 10'd109) & ~(trunc_ln321_fu_7683_p1 == 10'd108) & ~(trunc_ln321_fu_7683_p1 == 10'd107) & ~(trunc_ln321_fu_7683_p1 == 10'd106) & ~(trunc_ln321_fu_7683_p1 == 10'd105) & ~(trunc_ln321_fu_7683_p1 == 10'd104) & ~(trunc_ln321_fu_7683_p1 == 10'd103) & ~(trunc_ln321_fu_7683_p1 == 10'd102) & ~(trunc_ln321_fu_7683_p1 == 10'd101) & ~(trunc_ln321_fu_7683_p1 == 10'd100) & ~(trunc_ln321_fu_7683_p1 == 10'd99) & ~(trunc_ln321_fu_7683_p1 == 10'd98) & ~(trunc_ln321_fu_7683_p1 == 10'd97) & ~(trunc_ln321_fu_7683_p1 == 10'd96) & ~(trunc_ln321_fu_7683_p1 == 10'd95) & ~(trunc_ln321_fu_7683_p1 == 10'd94) & ~(trunc_ln321_fu_7683_p1 == 10'd93) & ~(trunc_ln321_fu_7683_p1 == 10'd92) & ~(trunc_ln321_fu_7683_p1 == 10'd91) & ~(trunc_ln321_fu_7683_p1 == 10'd90) & ~(trunc_ln321_fu_7683_p1 == 10'd89) & ~(trunc_ln321_fu_7683_p1 == 10'd88) & ~(trunc_ln321_fu_7683_p1 == 10'd87) & ~(trunc_ln321_fu_7683_p1 == 10'd86) & ~(trunc_ln321_fu_7683_p1 == 10'd85) & ~(trunc_ln321_fu_7683_p1 == 10'd84) & ~(trunc_ln321_fu_7683_p1 == 10'd83) & ~(trunc_ln321_fu_7683_p1 == 10'd82) & ~(trunc_ln321_fu_7683_p1 == 10'd81) & ~(trunc_ln321_fu_7683_p1 == 10'd80) & ~(trunc_ln321_fu_7683_p1 == 10'd79) & ~(trunc_ln321_fu_7683_p1 == 10'd78) & ~(trunc_ln321_fu_7683_p1 == 10'd77) & ~(trunc_ln321_fu_7683_p1 == 10'd76) & ~(trunc_ln321_fu_7683_p1 == 10'd75) & ~(trunc_ln321_fu_7683_p1 == 10'd74) & ~(trunc_ln321_fu_7683_p1 == 10'd73) & ~(trunc_ln321_fu_7683_p1 == 10'd72) & ~(trunc_ln321_fu_7683_p1 == 10'd71) & ~(trunc_ln321_fu_7683_p1 == 10'd70) & ~(trunc_ln321_fu_7683_p1 == 10'd69) & ~(trunc_ln321_fu_7683_p1 == 10'd68) & ~(trunc_ln321_fu_7683_p1 == 10'd67) & ~(trunc_ln321_fu_7683_p1 == 10'd66) & ~(trunc_ln321_fu_7683_p1 == 10'd65) & ~(trunc_ln321_fu_7683_p1 == 10'd64) & ~(trunc_ln321_fu_7683_p1 == 10'd63) & ~(trunc_ln321_fu_7683_p1 == 10'd62) & ~(trunc_ln321_fu_7683_p1 == 10'd61) & ~(trunc_ln321_fu_7683_p1 == 10'd60) & ~(trunc_ln321_fu_7683_p1 == 10'd59) & ~(trunc_ln321_fu_7683_p1 == 10'd58) & ~(trunc_ln321_fu_7683_p1 == 10'd57) & ~(trunc_ln321_fu_7683_p1 == 10'd56) & ~(trunc_ln321_fu_7683_p1 == 10'd55) & ~(trunc_ln321_fu_7683_p1 == 10'd54) & ~(trunc_ln321_fu_7683_p1 == 10'd53) & ~(trunc_ln321_fu_7683_p1 == 10'd52) & ~(trunc_ln321_fu_7683_p1 == 10'd51) & ~(trunc_ln321_fu_7683_p1 == 10'd50) & ~(trunc_ln321_fu_7683_p1 == 10'd49) & ~(trunc_ln321_fu_7683_p1 == 10'd48) & ~(trunc_ln321_fu_7683_p1 == 10'd47) & ~(trunc_ln321_fu_7683_p1 == 10'd46) & ~(trunc_ln321_fu_7683_p1 == 10'd45) & ~(trunc_ln321_fu_7683_p1 == 10'd44) & ~(trunc_ln321_fu_7683_p1 == 10'd43) & ~(trunc_ln321_fu_7683_p1 == 10'd42) & ~(trunc_ln321_fu_7683_p1 == 10'd41) & ~(trunc_ln321_fu_7683_p1 == 10'd40) & ~(trunc_ln321_fu_7683_p1 == 10'd39) & ~(trunc_ln321_fu_7683_p1 == 10'd38) & ~(trunc_ln321_fu_7683_p1 == 10'd37) & ~(trunc_ln321_fu_7683_p1 == 10'd36) & ~(trunc_ln321_fu_7683_p1 == 10'd35) & ~(trunc_ln321_fu_7683_p1 == 10'd34) & ~(trunc_ln321_fu_7683_p1 == 10'd33) & ~(trunc_ln321_fu_7683_p1 == 10'd32) & ~(trunc_ln321_fu_7683_p1 == 10'd31) & ~(trunc_ln321_fu_7683_p1 == 10'd30) & ~(trunc_ln321_fu_7683_p1 == 10'd29) & ~(trunc_ln321_fu_7683_p1 == 10'd28) & ~(trunc_ln321_fu_7683_p1 == 10'd27) & ~(trunc_ln321_fu_7683_p1 == 10'd26) & ~(trunc_ln321_fu_7683_p1 == 10'd574) & ~(trunc_ln321_fu_7683_p1 == 10'd573) & ~(trunc_ln321_fu_7683_p1 == 10'd572) & ~(trunc_ln321_fu_7683_p1 == 10'd25) & ~(trunc_ln321_fu_7683_p1 == 10'd571) & ~(trunc_ln321_fu_7683_p1 == 10'd570) & ~(trunc_ln321_fu_7683_p1 == 10'd569) & ~(trunc_ln321_fu_7683_p1 == 10'd568) & ~(trunc_ln321_fu_7683_p1 == 10'd567) & ~(trunc_ln321_fu_7683_p1 == 10'd566) & ~(trunc_ln321_fu_7683_p1 == 10'd565) & ~(trunc_ln321_fu_7683_p1 == 10'd564) & ~(trunc_ln321_fu_7683_p1 == 10'd563) & ~(trunc_ln321_fu_7683_p1 == 10'd562) & ~(trunc_ln321_fu_7683_p1 == 10'd24) & ~(trunc_ln321_fu_7683_p1 == 10'd561) & ~(trunc_ln321_fu_7683_p1 == 10'd560) & ~(trunc_ln321_fu_7683_p1 == 10'd559) & ~(trunc_ln321_fu_7683_p1 == 10'd558) & ~(trunc_ln321_fu_7683_p1 == 10'd557) & ~(trunc_ln321_fu_7683_p1 == 10'd556) & ~(trunc_ln321_fu_7683_p1 == 10'd555) & ~(trunc_ln321_fu_7683_p1 == 10'd554) & ~(trunc_ln321_fu_7683_p1 == 10'd553) & ~(trunc_ln321_fu_7683_p1 == 10'd552) & ~(trunc_ln321_fu_7683_p1 == 10'd23) & ~(trunc_ln321_fu_7683_p1 == 10'd551) & ~(trunc_ln321_fu_7683_p1 == 10'd550) & ~(trunc_ln321_fu_7683_p1 == 10'd549) & ~(trunc_ln321_fu_7683_p1 == 10'd548) & ~(trunc_ln321_fu_7683_p1 == 10'd547) & ~(trunc_ln321_fu_7683_p1 == 10'd546) & ~(trunc_ln321_fu_7683_p1 == 10'd545) & ~(trunc_ln321_fu_7683_p1 == 10'd544) & ~(trunc_ln321_fu_7683_p1 == 10'd543) & ~(trunc_ln321_fu_7683_p1 == 10'd542) & ~(trunc_ln321_fu_7683_p1 == 10'd22) & ~(trunc_ln321_fu_7683_p1 == 10'd541) & ~(trunc_ln321_fu_7683_p1 == 10'd540) & ~(trunc_ln321_fu_7683_p1 == 10'd539) & ~(trunc_ln321_fu_7683_p1 == 10'd538) & ~(trunc_ln321_fu_7683_p1 == 10'd537) & ~(trunc_ln321_fu_7683_p1 == 10'd536) & ~(trunc_ln321_fu_7683_p1 == 10'd535) & ~(trunc_ln321_fu_7683_p1 == 10'd534) & ~(trunc_ln321_fu_7683_p1 == 10'd533) & ~(trunc_ln321_fu_7683_p1 == 10'd532) & ~(trunc_ln321_fu_7683_p1 == 10'd21) & ~(trunc_ln321_fu_7683_p1 == 10'd531) & ~(trunc_ln321_fu_7683_p1 == 10'd530) & ~(trunc_ln321_fu_7683_p1 == 10'd529) & ~(trunc_ln321_fu_7683_p1 == 10'd528) & ~(trunc_ln321_fu_7683_p1 == 10'd527) & ~(trunc_ln321_fu_7683_p1 == 10'd526) & ~(trunc_ln321_fu_7683_p1 == 10'd525) & ~(trunc_ln321_fu_7683_p1 == 10'd524) & ~(trunc_ln321_fu_7683_p1 == 10'd523) & ~(trunc_ln321_fu_7683_p1 == 10'd522) & ~(trunc_ln321_fu_7683_p1 == 10'd20) & ~(trunc_ln321_fu_7683_p1 == 10'd521) & ~(trunc_ln321_fu_7683_p1 == 10'd520) & ~(trunc_ln321_fu_7683_p1 == 10'd519) & ~(trunc_ln321_fu_7683_p1 == 10'd518) & ~(trunc_ln321_fu_7683_p1 == 10'd517) & ~(trunc_ln321_fu_7683_p1 == 10'd516) & ~(trunc_ln321_fu_7683_p1 == 10'd515) & ~(trunc_ln321_fu_7683_p1 == 10'd514) & ~(trunc_ln321_fu_7683_p1 == 10'd513) & ~(trunc_ln321_fu_7683_p1 == 10'd512) & ~(trunc_ln321_fu_7683_p1 == 10'd19) & ~(trunc_ln321_fu_7683_p1 == 10'd511) & ~(trunc_ln321_fu_7683_p1 == 10'd510) & ~(trunc_ln321_fu_7683_p1 == 10'd509) & ~(trunc_ln321_fu_7683_p1 == 10'd508) & ~(trunc_ln321_fu_7683_p1 == 10'd507) & ~(trunc_ln321_fu_7683_p1 == 10'd506) & ~(trunc_ln321_fu_7683_p1 == 10'd505) & ~(trunc_ln321_fu_7683_p1 == 10'd504) & ~(trunc_ln321_fu_7683_p1 == 10'd503) & ~(trunc_ln321_fu_7683_p1 == 10'd502) & ~(trunc_ln321_fu_7683_p1 == 10'd18) & ~(trunc_ln321_fu_7683_p1 == 10'd501) & ~(trunc_ln321_fu_7683_p1 == 10'd500) & ~(trunc_ln321_fu_7683_p1 == 10'd499) & ~(trunc_ln321_fu_7683_p1 == 10'd498) & ~(trunc_ln321_fu_7683_p1 == 10'd497) & ~(trunc_ln321_fu_7683_p1 == 10'd496) & ~(trunc_ln321_fu_7683_p1 == 10'd495) & ~(trunc_ln321_fu_7683_p1 == 10'd494) & ~(trunc_ln321_fu_7683_p1 == 10'd493) & ~(trunc_ln321_fu_7683_p1 == 10'd492) & ~(trunc_ln321_fu_7683_p1 == 10'd17) & ~(trunc_ln321_fu_7683_p1 == 10'd491) & ~(trunc_ln321_fu_7683_p1 == 10'd490) & ~(trunc_ln321_fu_7683_p1 == 10'd489) & ~(trunc_ln321_fu_7683_p1 == 10'd488) & ~(trunc_ln321_fu_7683_p1 == 10'd487) & ~(trunc_ln321_fu_7683_p1 == 10'd486) & ~(trunc_ln321_fu_7683_p1 == 10'd485) & ~(trunc_ln321_fu_7683_p1 == 10'd484) & ~(trunc_ln321_fu_7683_p1 == 10'd483) & ~(trunc_ln321_fu_7683_p1 == 10'd482) & ~(trunc_ln321_fu_7683_p1 == 10'd16) & ~(trunc_ln321_fu_7683_p1 == 10'd481) & ~(trunc_ln321_fu_7683_p1 == 10'd480) & ~(trunc_ln321_fu_7683_p1 == 10'd479) & ~(trunc_ln321_fu_7683_p1 == 10'd478) & ~(trunc_ln321_fu_7683_p1 == 10'd477) & ~(trunc_ln321_fu_7683_p1 == 10'd476) & ~(trunc_ln321_fu_7683_p1 == 10'd475) & ~(trunc_ln321_fu_7683_p1 == 10'd474) & ~(trunc_ln321_fu_7683_p1 == 10'd473) & ~(trunc_ln321_fu_7683_p1 == 10'd472) & ~(trunc_ln321_fu_7683_p1 == 10'd15) & ~(trunc_ln321_fu_7683_p1 == 10'd471) & ~(trunc_ln321_fu_7683_p1 == 10'd470) & ~(trunc_ln321_fu_7683_p1 == 10'd469) & ~(trunc_ln321_fu_7683_p1 == 10'd468) & ~(trunc_ln321_fu_7683_p1 == 10'd467) & ~(trunc_ln321_fu_7683_p1 == 10'd466) & ~(trunc_ln321_fu_7683_p1 == 10'd465) & ~(trunc_ln321_fu_7683_p1 == 10'd464) & ~(trunc_ln321_fu_7683_p1 == 10'd463) & ~(trunc_ln321_fu_7683_p1 == 10'd462) & ~(trunc_ln321_fu_7683_p1 == 10'd14) & ~(trunc_ln321_fu_7683_p1 == 10'd461) & ~(trunc_ln321_fu_7683_p1 == 10'd460) & ~(trunc_ln321_fu_7683_p1 == 10'd459) & ~(trunc_ln321_fu_7683_p1 == 10'd458) & ~(trunc_ln321_fu_7683_p1 == 10'd457) & ~(trunc_ln321_fu_7683_p1 == 10'd456) & ~(trunc_ln321_fu_7683_p1 == 10'd455) & ~(trunc_ln321_fu_7683_p1 == 10'd454) & ~(trunc_ln321_fu_7683_p1 == 10'd453) & ~(trunc_ln321_fu_7683_p1 == 10'd452) & ~(trunc_ln321_fu_7683_p1 == 10'd13) & ~(trunc_ln321_fu_7683_p1 == 10'd451) & ~(trunc_ln321_fu_7683_p1 == 10'd450) & ~(trunc_ln321_fu_7683_p1 == 10'd449) & ~(trunc_ln321_fu_7683_p1 == 10'd448) & ~(trunc_ln321_fu_7683_p1 == 10'd447) & ~(trunc_ln321_fu_7683_p1 == 10'd446) & ~(trunc_ln321_fu_7683_p1 == 10'd445) & ~(trunc_ln321_fu_7683_p1 == 10'd444) & ~(trunc_ln321_fu_7683_p1 == 10'd443) & ~(trunc_ln321_fu_7683_p1 == 10'd442) & ~(trunc_ln321_fu_7683_p1 == 10'd12) & ~(trunc_ln321_fu_7683_p1 == 10'd441) & ~(trunc_ln321_fu_7683_p1 == 10'd440) & ~(trunc_ln321_fu_7683_p1 == 10'd439) & ~(trunc_ln321_fu_7683_p1 == 10'd438) & ~(trunc_ln321_fu_7683_p1 == 10'd437) & ~(trunc_ln321_fu_7683_p1 == 10'd436) & ~(trunc_ln321_fu_7683_p1 == 10'd435) & ~(trunc_ln321_fu_7683_p1 == 10'd434) & ~(trunc_ln321_fu_7683_p1 == 10'd433) & ~(trunc_ln321_fu_7683_p1 == 10'd432) & ~(trunc_ln321_fu_7683_p1 == 10'd11) & ~(trunc_ln321_fu_7683_p1 == 10'd431) & ~(trunc_ln321_fu_7683_p1 == 10'd430) & ~(trunc_ln321_fu_7683_p1 == 10'd429) & ~(trunc_ln321_fu_7683_p1 == 10'd428) & ~(trunc_ln321_fu_7683_p1 == 10'd427) & ~(trunc_ln321_fu_7683_p1 == 10'd426) & ~(trunc_ln321_fu_7683_p1 == 10'd425) & ~(trunc_ln321_fu_7683_p1 == 10'd424) & ~(trunc_ln321_fu_7683_p1 == 10'd423) & ~(trunc_ln321_fu_7683_p1 == 10'd422) & ~(trunc_ln321_fu_7683_p1 == 10'd10) & ~(trunc_ln321_fu_7683_p1 == 10'd421) & ~(trunc_ln321_fu_7683_p1 == 10'd420) & ~(trunc_ln321_fu_7683_p1 == 10'd419) & ~(trunc_ln321_fu_7683_p1 == 10'd418) & ~(trunc_ln321_fu_7683_p1 == 10'd417) & ~(trunc_ln321_fu_7683_p1 == 10'd416) & ~(trunc_ln321_fu_7683_p1 == 10'd415) & ~(trunc_ln321_fu_7683_p1 == 10'd414) & ~(trunc_ln321_fu_7683_p1 == 10'd413) & ~(trunc_ln321_fu_7683_p1 == 10'd412) & ~(trunc_ln321_fu_7683_p1 == 10'd9) & ~(trunc_ln321_fu_7683_p1 == 10'd411) & ~(trunc_ln321_fu_7683_p1 == 10'd410) & ~(trunc_ln321_fu_7683_p1 == 10'd409) & ~(trunc_ln321_fu_7683_p1 == 10'd408) & ~(trunc_ln321_fu_7683_p1 == 10'd407) & ~(trunc_ln321_fu_7683_p1 == 10'd406) & ~(trunc_ln321_fu_7683_p1 == 10'd405) & ~(trunc_ln321_fu_7683_p1 == 10'd404) & ~(trunc_ln321_fu_7683_p1 == 10'd403) & ~(trunc_ln321_fu_7683_p1 == 10'd402) & ~(trunc_ln321_fu_7683_p1 == 10'd8) & ~(trunc_ln321_fu_7683_p1 == 10'd401) & ~(trunc_ln321_fu_7683_p1 == 10'd400) & ~(trunc_ln321_fu_7683_p1 == 10'd399) & ~(trunc_ln321_fu_7683_p1 == 10'd398) & ~(trunc_ln321_fu_7683_p1 == 10'd397) & ~(trunc_ln321_fu_7683_p1 == 10'd396) & ~(trunc_ln321_fu_7683_p1 == 10'd395) & ~(trunc_ln321_fu_7683_p1 == 10'd394) & ~(trunc_ln321_fu_7683_p1 == 10'd393) & ~(trunc_ln321_fu_7683_p1 == 10'd392) & ~(trunc_ln321_fu_7683_p1 == 10'd7) & ~(trunc_ln321_fu_7683_p1 == 10'd391) & ~(trunc_ln321_fu_7683_p1 == 10'd390) & ~(trunc_ln321_fu_7683_p1 == 10'd389) & ~(trunc_ln321_fu_7683_p1 == 10'd388) & ~(trunc_ln321_fu_7683_p1 == 10'd387) & ~(trunc_ln321_fu_7683_p1 == 10'd386) & ~(trunc_ln321_fu_7683_p1 == 10'd385) & ~(trunc_ln321_fu_7683_p1 == 10'd384) & ~(trunc_ln321_fu_7683_p1 == 10'd383) & ~(trunc_ln321_fu_7683_p1 == 10'd382) & ~(trunc_ln321_fu_7683_p1 == 10'd6) & ~(trunc_ln321_fu_7683_p1 == 10'd381) & ~(trunc_ln321_fu_7683_p1 == 10'd380) & ~(trunc_ln321_fu_7683_p1 == 10'd379) & ~(trunc_ln321_fu_7683_p1 == 10'd378) & ~(trunc_ln321_fu_7683_p1 == 10'd377) & ~(trunc_ln321_fu_7683_p1 == 10'd376) & ~(trunc_ln321_fu_7683_p1 == 10'd375) & ~(trunc_ln321_fu_7683_p1 == 10'd374) & ~(trunc_ln321_fu_7683_p1 == 10'd373) & ~(trunc_ln321_fu_7683_p1 == 10'd372) & ~(trunc_ln321_fu_7683_p1 == 10'd5) & ~(trunc_ln321_fu_7683_p1 == 10'd371) & ~(trunc_ln321_fu_7683_p1 == 10'd370) & ~(trunc_ln321_fu_7683_p1 == 10'd369) & ~(trunc_ln321_fu_7683_p1 == 10'd368) & ~(trunc_ln321_fu_7683_p1 == 10'd367) & ~(trunc_ln321_fu_7683_p1 == 10'd366) & ~(trunc_ln321_fu_7683_p1 == 10'd365) & ~(trunc_ln321_fu_7683_p1 == 10'd364) & ~(trunc_ln321_fu_7683_p1 == 10'd363) & ~(trunc_ln321_fu_7683_p1 == 10'd362) & ~(trunc_ln321_fu_7683_p1 == 10'd4) & ~(trunc_ln321_fu_7683_p1 == 10'd361) & ~(trunc_ln321_fu_7683_p1 == 10'd360) & ~(trunc_ln321_fu_7683_p1 == 10'd359) & ~(trunc_ln321_fu_7683_p1 == 10'd358) & ~(trunc_ln321_fu_7683_p1 == 10'd357) & ~(trunc_ln321_fu_7683_p1 == 10'd356) & ~(trunc_ln321_fu_7683_p1 == 10'd355) & ~(trunc_ln321_fu_7683_p1 == 10'd354) & ~(trunc_ln321_fu_7683_p1 == 10'd353) & ~(trunc_ln321_fu_7683_p1 == 10'd352) & ~(trunc_ln321_fu_7683_p1 == 10'd3) & ~(trunc_ln321_fu_7683_p1 == 10'd351) & ~(trunc_ln321_fu_7683_p1 == 10'd350) & ~(trunc_ln321_fu_7683_p1 == 10'd349) & ~(trunc_ln321_fu_7683_p1 == 10'd348) & ~(trunc_ln321_fu_7683_p1 == 10'd347) & ~(trunc_ln321_fu_7683_p1 == 10'd346) & ~(trunc_ln321_fu_7683_p1 == 10'd345) & ~(trunc_ln321_fu_7683_p1 == 10'd344) & ~(trunc_ln321_fu_7683_p1 == 10'd343) & ~(trunc_ln321_fu_7683_p1 == 10'd342) & ~(trunc_ln321_fu_7683_p1 == 10'd2) & ~(trunc_ln321_fu_7683_p1 == 10'd341) & ~(trunc_ln321_fu_7683_p1 == 10'd340) & ~(trunc_ln321_fu_7683_p1 == 10'd339) & ~(trunc_ln321_fu_7683_p1 == 10'd338) & ~(trunc_ln321_fu_7683_p1 == 10'd337) & ~(trunc_ln321_fu_7683_p1 == 10'd336) & ~(trunc_ln321_fu_7683_p1 == 10'd335) & ~(trunc_ln321_fu_7683_p1 == 10'd334) & ~(trunc_ln321_fu_7683_p1 == 10'd333) & ~(trunc_ln321_fu_7683_p1 == 10'd332) & ~(trunc_ln321_fu_7683_p1 == 10'd1) & ~(trunc_ln321_fu_7683_p1 == 10'd331) & ~(trunc_ln321_fu_7683_p1 == 10'd330) & ~(trunc_ln321_fu_7683_p1 == 10'd329) & ~(trunc_ln321_fu_7683_p1 == 10'd328) & ~(trunc_ln321_fu_7683_p1 == 10'd327) & ~(trunc_ln321_fu_7683_p1 == 10'd326) & ~(trunc_ln321_fu_7683_p1 == 10'd325) & ~(trunc_ln321_fu_7683_p1 == 10'd324) & ~(trunc_ln321_fu_7683_p1 == 10'd323) & ~(trunc_ln321_fu_7683_p1 == 10'd322) & ~(trunc_ln321_fu_7683_p1 == 10'd0) & ~(trunc_ln321_fu_7683_p1 == 10'd321) & ~(trunc_ln321_fu_7683_p1 == 10'd320) & ~(trunc_ln321_fu_7683_p1 == 10'd319) & ~(trunc_ln321_fu_7683_p1 == 10'd318) & ~(trunc_ln321_fu_7683_p1 == 10'd317) & ~(trunc_ln321_fu_7683_p1 == 10'd316) & ~(trunc_ln321_fu_7683_p1 == 10'd315) & ~(trunc_ln321_fu_7683_p1 == 10'd314) & ~(trunc_ln321_fu_7683_p1 == 10'd313) & ~(trunc_ln321_fu_7683_p1 == 10'd312) & ~(trunc_ln321_fu_7683_p1 == 10'd311) & ~(trunc_ln321_fu_7683_p1 == 10'd310) & ~(trunc_ln321_fu_7683_p1 == 10'd309) & ~(trunc_ln321_fu_7683_p1 == 10'd308) & ~(trunc_ln321_fu_7683_p1 == 10'd307) & ~(trunc_ln321_fu_7683_p1 == 10'd306) & ~(trunc_ln321_fu_7683_p1 == 10'd305) & ~(trunc_ln321_fu_7683_p1 == 10'd304) & ~(trunc_ln321_fu_7683_p1 == 10'd303) & ~(trunc_ln321_fu_7683_p1 == 10'd302) & ~(trunc_ln321_fu_7683_p1 == 10'd301) & ~(trunc_ln321_fu_7683_p1 == 10'd300) & ~(trunc_ln321_fu_7683_p1 == 10'd299) & ~(trunc_ln321_fu_7683_p1 == 10'd298) & ~(trunc_ln321_fu_7683_p1 == 10'd297) & ~(trunc_ln321_fu_7683_p1 == 10'd296) & ~(trunc_ln321_fu_7683_p1 == 10'd295) & ~(trunc_ln321_fu_7683_p1 == 10'd294) & ~(trunc_ln321_fu_7683_p1 == 10'd293) & ~(trunc_ln321_fu_7683_p1 == 10'd292) & ~(trunc_ln321_fu_7683_p1 == 10'd291) & ~(trunc_ln321_fu_7683_p1 == 10'd290) & ~(trunc_ln321_fu_7683_p1 == 10'd289) & ~(trunc_ln321_fu_7683_p1 == 10'd288) & ~(trunc_ln321_fu_7683_p1 == 10'd287) & ~(trunc_ln321_fu_7683_p1 == 10'd286) & ~(trunc_ln321_fu_7683_p1 == 10'd285) & ~(trunc_ln321_fu_7683_p1 == 10'd284) & ~(trunc_ln321_fu_7683_p1 == 10'd283) & ~(trunc_ln321_fu_7683_p1 == 10'd282) & ~(trunc_ln321_fu_7683_p1 == 10'd281) & ~(trunc_ln321_fu_7683_p1 == 10'd280) & ~(trunc_ln321_fu_7683_p1 == 10'd279) & ~(trunc_ln321_fu_7683_p1 == 10'd278) & ~(trunc_ln321_fu_7683_p1 == 10'd277) & ~(trunc_ln321_fu_7683_p1 == 10'd276) & ~(trunc_ln321_fu_7683_p1 == 10'd275) & ~(trunc_ln321_fu_7683_p1 == 10'd274) & ~(trunc_ln321_fu_7683_p1 == 10'd273) & ~(trunc_ln321_fu_7683_p1 == 10'd272) & ~(trunc_ln321_fu_7683_p1 == 10'd271) & ~(trunc_ln321_fu_7683_p1 == 10'd270) & ~(trunc_ln321_fu_7683_p1 == 10'd269) & ~(trunc_ln321_fu_7683_p1 == 10'd268) & ~(trunc_ln321_fu_7683_p1 == 10'd267) & ~(trunc_ln321_fu_7683_p1 == 10'd266) & ~(trunc_ln321_fu_7683_p1 == 10'd265) & ~(trunc_ln321_fu_7683_p1 == 10'd264) & ~(trunc_ln321_fu_7683_p1 == 10'd263) & ~(trunc_ln321_fu_7683_p1 == 10'd262) & ~(trunc_ln321_fu_7683_p1 == 10'd261) & ~(trunc_ln321_fu_7683_p1 == 10'd260) & ~(trunc_ln321_fu_7683_p1 == 10'd259) & ~(trunc_ln321_fu_7683_p1 == 10'd258) & ~(trunc_ln321_fu_7683_p1 == 10'd257) & ~(trunc_ln321_fu_7683_p1 == 10'd256) & ~(trunc_ln321_fu_7683_p1 == 10'd255) & ~(trunc_ln321_fu_7683_p1 == 10'd254) & ~(trunc_ln321_fu_7683_p1 == 10'd253) & ~(trunc_ln321_fu_7683_p1 == 10'd252) & ~(trunc_ln321_fu_7683_p1 == 10'd251) & ~(trunc_ln321_fu_7683_p1 == 10'd250) & ~(trunc_ln321_fu_7683_p1 == 10'd249) & ~(trunc_ln321_fu_7683_p1 == 10'd248) & ~(trunc_ln321_fu_7683_p1 == 10'd247) & ~(trunc_ln321_fu_7683_p1 == 10'd246) & ~(trunc_ln321_fu_7683_p1 == 10'd245) & ~(trunc_ln321_fu_7683_p1 == 10'd244) & ~(trunc_ln321_fu_7683_p1 == 10'd243) & ~(trunc_ln321_fu_7683_p1 == 10'd242) & ~(trunc_ln321_fu_7683_p1 == 10'd241) & ~(trunc_ln321_fu_7683_p1 == 10'd240) & ~(trunc_ln321_fu_7683_p1 == 10'd239) & ~(trunc_ln321_fu_7683_p1 == 10'd238) & ~(trunc_ln321_fu_7683_p1 == 10'd237) & ~(trunc_ln321_fu_7683_p1 == 10'd236) & ~(trunc_ln321_fu_7683_p1 == 10'd235) & ~(trunc_ln321_fu_7683_p1 == 10'd234) & ~(trunc_ln321_fu_7683_p1 == 10'd233) & ~(trunc_ln321_fu_7683_p1 == 10'd232) & ~(trunc_ln321_fu_7683_p1 == 10'd231) & ~(trunc_ln321_fu_7683_p1 == 10'd230) & ~(trunc_ln321_fu_7683_p1 == 10'd229) & ~(trunc_ln321_fu_7683_p1 == 10'd228) & ~(trunc_ln321_fu_7683_p1 == 10'd227) & ~(trunc_ln321_fu_7683_p1 == 10'd226) & ~(trunc_ln321_fu_7683_p1 == 10'd225) & ~(trunc_ln321_fu_7683_p1 == 10'd224) & ~(trunc_ln321_fu_7683_p1 == 10'd223) & ~(trunc_ln321_fu_7683_p1 == 10'd222) & ~(trunc_ln321_fu_7683_p1 == 10'd221) & ~(trunc_ln321_fu_7683_p1 == 10'd220) & ~(trunc_ln321_fu_7683_p1 == 10'd219) & ~(trunc_ln321_fu_7683_p1 == 10'd218) & ~(trunc_ln321_fu_7683_p1 == 10'd217) & ~(trunc_ln321_fu_7683_p1 == 10'd216) & ~(trunc_ln321_fu_7683_p1 == 10'd215) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd326)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd325)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd324)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd323)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd322)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd321)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd320)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd319)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd318)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd317)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd316)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd315)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd314)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd313)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd312)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd311)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd310)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd309)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd308)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd307)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd306)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd305)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd304)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd303)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd302)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd301)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd300)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd299)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd298)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd297)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd296)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd295)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd294)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd293)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd292)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd291)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd290)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd289)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd288)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd287)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd286)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd285)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd284)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd283)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd282)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd281)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd280)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd279)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd278)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd277)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd276)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd275)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd274)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd273)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd272)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd271)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd270)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd269)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd268)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd267)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd266)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd265)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd264)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd263)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd262)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd261)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd260)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd259)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd258)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd257)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd256)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd255)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd254)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd253)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd252)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd251)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd250)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd249)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd248)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd247)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd246)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd245)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd244)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd243)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd242)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd241)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd240)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd239)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd238)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd237)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd236)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd235)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd234)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd233)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd232)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd231)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd230)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd229)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd228)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd227)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd226)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd225)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd224)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd223)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd222)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd221)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd220)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd219)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd218)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd217)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd216)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd215)))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_3600 <= in_V_V_TDATA;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_3600 <= ap_phi_reg_pp0_iter0_act_m_val_V_reg_3600;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_reg_3589 <= i_fu_4775_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_reg_3589 <= 21'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_15104 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        nf_0_fu_3566 <= select_ln301_fu_10945_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        nf_0_fu_3566 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_10656_p2 == 1'd0) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        sf_1_fu_1258 <= sf_fu_10650_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_10656_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        sf_1_fu_1258 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        accu_0_0_V_1_fu_1242 <= accu_0_0_V_fu_10765_p2;
        accu_0_1_V_1_fu_1246 <= accu_0_1_V_fu_10807_p2;
        accu_0_2_V_1_fu_1250 <= accu_0_2_V_fu_10849_p2;
        accu_0_3_V_1_fu_1254 <= accu_0_3_V_fu_10891_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_4769_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln271_reg_15056 <= icmp_ln271_fu_10570_p2;
        icmp_ln289_reg_15104 <= icmp_ln289_fu_10656_p2;
        p_Result_1_0_1_reg_15069 <= {{weight_V_V_TDATA[7:4]}};
        p_Result_1_1_1_reg_15079 <= {{weight_V_V_TDATA[15:12]}};
        p_Result_1_1_reg_15074 <= {{weight_V_V_TDATA[11:8]}};
        p_Result_1_2_1_reg_15089 <= {{weight_V_V_TDATA[23:20]}};
        p_Result_1_2_reg_15084 <= {{weight_V_V_TDATA[19:16]}};
        p_Result_1_3_1_reg_15099 <= {{weight_V_V_TDATA[31:28]}};
        p_Result_1_3_reg_15094 <= {{weight_V_V_TDATA[27:24]}};
        trunc_ln647_reg_15064 <= trunc_ln647_fu_10576_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd99))) begin
        tmp_V_100_fu_1658 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd100))) begin
        tmp_V_101_fu_1662 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd101))) begin
        tmp_V_102_fu_1666 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd102))) begin
        tmp_V_103_fu_1670 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd103))) begin
        tmp_V_104_fu_1674 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd104))) begin
        tmp_V_105_fu_1678 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd105))) begin
        tmp_V_106_fu_1682 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd106))) begin
        tmp_V_107_fu_1686 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd107))) begin
        tmp_V_108_fu_1690 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd108))) begin
        tmp_V_109_fu_1694 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd9))) begin
        tmp_V_10_fu_1298 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd109))) begin
        tmp_V_110_fu_1698 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd110))) begin
        tmp_V_111_fu_1702 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd111))) begin
        tmp_V_112_fu_1706 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd112))) begin
        tmp_V_113_fu_1710 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd113))) begin
        tmp_V_114_fu_1714 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd114))) begin
        tmp_V_115_fu_1718 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd115))) begin
        tmp_V_116_fu_1722 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd116))) begin
        tmp_V_117_fu_1726 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd117))) begin
        tmp_V_118_fu_1730 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd118))) begin
        tmp_V_119_fu_1734 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd10))) begin
        tmp_V_11_fu_1302 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd119))) begin
        tmp_V_120_fu_1738 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd120))) begin
        tmp_V_121_fu_1742 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd121))) begin
        tmp_V_122_fu_1746 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd122))) begin
        tmp_V_123_fu_1750 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd123))) begin
        tmp_V_124_fu_1754 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd124))) begin
        tmp_V_125_fu_1758 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd125))) begin
        tmp_V_126_fu_1762 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd126))) begin
        tmp_V_127_fu_1766 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd127))) begin
        tmp_V_128_fu_1770 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd128))) begin
        tmp_V_129_fu_1774 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd11))) begin
        tmp_V_12_fu_1306 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd129))) begin
        tmp_V_130_fu_1778 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd130))) begin
        tmp_V_131_fu_1782 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd131))) begin
        tmp_V_132_fu_1786 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd132))) begin
        tmp_V_133_fu_1790 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd133))) begin
        tmp_V_134_fu_1794 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd134))) begin
        tmp_V_135_fu_1798 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd135))) begin
        tmp_V_136_fu_1802 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd136))) begin
        tmp_V_137_fu_1806 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd137))) begin
        tmp_V_138_fu_1810 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd138))) begin
        tmp_V_139_fu_1814 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd12))) begin
        tmp_V_13_fu_1310 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd139))) begin
        tmp_V_140_fu_1818 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd140))) begin
        tmp_V_141_fu_1822 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd141))) begin
        tmp_V_142_fu_1826 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd142))) begin
        tmp_V_143_fu_1830 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd143))) begin
        tmp_V_144_fu_1834 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd144))) begin
        tmp_V_145_fu_1838 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd145))) begin
        tmp_V_146_fu_1842 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd146))) begin
        tmp_V_147_fu_1846 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd147))) begin
        tmp_V_148_fu_1850 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd148))) begin
        tmp_V_149_fu_1854 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd13))) begin
        tmp_V_14_fu_1314 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd149))) begin
        tmp_V_150_fu_1858 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd150))) begin
        tmp_V_151_fu_1862 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd151))) begin
        tmp_V_152_fu_1866 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd152))) begin
        tmp_V_153_fu_1870 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd153))) begin
        tmp_V_154_fu_1874 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd154))) begin
        tmp_V_155_fu_1878 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd155))) begin
        tmp_V_156_fu_1882 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd156))) begin
        tmp_V_157_fu_1886 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd157))) begin
        tmp_V_158_fu_1890 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd158))) begin
        tmp_V_159_fu_1894 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd14))) begin
        tmp_V_15_fu_1318 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd159))) begin
        tmp_V_160_fu_1898 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd160))) begin
        tmp_V_161_fu_1902 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd161))) begin
        tmp_V_162_fu_1906 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd162))) begin
        tmp_V_163_fu_1910 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd163))) begin
        tmp_V_164_fu_1914 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd164))) begin
        tmp_V_165_fu_1918 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd165))) begin
        tmp_V_166_fu_1922 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd166))) begin
        tmp_V_167_fu_1926 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd167))) begin
        tmp_V_168_fu_1930 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd168))) begin
        tmp_V_169_fu_1934 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd15))) begin
        tmp_V_16_fu_1322 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd169))) begin
        tmp_V_170_fu_1938 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd170))) begin
        tmp_V_171_fu_1942 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd171))) begin
        tmp_V_172_fu_1946 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd172))) begin
        tmp_V_173_fu_1950 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd173))) begin
        tmp_V_174_fu_1954 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd174))) begin
        tmp_V_175_fu_1958 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd175))) begin
        tmp_V_176_fu_1962 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd176))) begin
        tmp_V_177_fu_1966 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd177))) begin
        tmp_V_178_fu_1970 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd178))) begin
        tmp_V_179_fu_1974 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd16))) begin
        tmp_V_17_fu_1326 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd179))) begin
        tmp_V_180_fu_1978 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd180))) begin
        tmp_V_181_fu_1982 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd181))) begin
        tmp_V_182_fu_1986 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd182))) begin
        tmp_V_183_fu_1990 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd183))) begin
        tmp_V_184_fu_1994 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd184))) begin
        tmp_V_185_fu_1998 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd185))) begin
        tmp_V_186_fu_2002 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd186))) begin
        tmp_V_187_fu_2006 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd187))) begin
        tmp_V_188_fu_2010 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd188))) begin
        tmp_V_189_fu_2014 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd17))) begin
        tmp_V_18_fu_1330 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd189))) begin
        tmp_V_190_fu_2018 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd190))) begin
        tmp_V_191_fu_2022 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd191))) begin
        tmp_V_192_fu_2026 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd192))) begin
        tmp_V_193_fu_2030 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd193))) begin
        tmp_V_194_fu_2034 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd194))) begin
        tmp_V_195_fu_2038 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd195))) begin
        tmp_V_196_fu_2042 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd196))) begin
        tmp_V_197_fu_2046 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd197))) begin
        tmp_V_198_fu_2050 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd198))) begin
        tmp_V_199_fu_2054 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd18))) begin
        tmp_V_19_fu_1334 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd1))) begin
        tmp_V_1_fu_1266 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd199))) begin
        tmp_V_200_fu_2058 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd200))) begin
        tmp_V_201_fu_2062 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd201))) begin
        tmp_V_202_fu_2066 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd202))) begin
        tmp_V_203_fu_2070 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd203))) begin
        tmp_V_204_fu_2074 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd204))) begin
        tmp_V_205_fu_2078 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd205))) begin
        tmp_V_206_fu_2082 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd206))) begin
        tmp_V_207_fu_2086 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd207))) begin
        tmp_V_208_fu_2090 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd208))) begin
        tmp_V_209_fu_2094 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd19))) begin
        tmp_V_20_fu_1338 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd209))) begin
        tmp_V_210_fu_2098 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd210))) begin
        tmp_V_211_fu_2102 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd211))) begin
        tmp_V_212_fu_2106 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd212))) begin
        tmp_V_213_fu_2110 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd213))) begin
        tmp_V_214_fu_2114 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd214))) begin
        tmp_V_215_fu_2118 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd215))) begin
        tmp_V_216_fu_2122 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd216))) begin
        tmp_V_217_fu_2126 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd217))) begin
        tmp_V_218_fu_2130 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd218))) begin
        tmp_V_219_fu_2134 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd20))) begin
        tmp_V_21_fu_1342 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd219))) begin
        tmp_V_220_fu_2138 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd220))) begin
        tmp_V_221_fu_2142 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd221))) begin
        tmp_V_222_fu_2146 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd222))) begin
        tmp_V_223_fu_2150 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd223))) begin
        tmp_V_224_fu_2154 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd224))) begin
        tmp_V_225_fu_2158 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd225))) begin
        tmp_V_226_fu_2162 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd226))) begin
        tmp_V_227_fu_2166 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd227))) begin
        tmp_V_228_fu_2170 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd228))) begin
        tmp_V_229_fu_2174 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd21))) begin
        tmp_V_22_fu_1346 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd229))) begin
        tmp_V_230_fu_2178 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd230))) begin
        tmp_V_231_fu_2182 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd231))) begin
        tmp_V_232_fu_2186 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd232))) begin
        tmp_V_233_fu_2190 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd233))) begin
        tmp_V_234_fu_2194 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd234))) begin
        tmp_V_235_fu_2198 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd235))) begin
        tmp_V_236_fu_2202 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd236))) begin
        tmp_V_237_fu_2206 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd237))) begin
        tmp_V_238_fu_2210 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd238))) begin
        tmp_V_239_fu_2214 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd22))) begin
        tmp_V_23_fu_1350 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd239))) begin
        tmp_V_240_fu_2218 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd240))) begin
        tmp_V_241_fu_2222 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd241))) begin
        tmp_V_242_fu_2226 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd242))) begin
        tmp_V_243_fu_2230 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd243))) begin
        tmp_V_244_fu_2234 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd244))) begin
        tmp_V_245_fu_2238 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd245))) begin
        tmp_V_246_fu_2242 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd246))) begin
        tmp_V_247_fu_2246 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd247))) begin
        tmp_V_248_fu_2250 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd248))) begin
        tmp_V_249_fu_2254 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd23))) begin
        tmp_V_24_fu_1354 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd249))) begin
        tmp_V_250_fu_2258 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd250))) begin
        tmp_V_251_fu_2262 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd251))) begin
        tmp_V_252_fu_2266 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd252))) begin
        tmp_V_253_fu_2270 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd253))) begin
        tmp_V_254_fu_2274 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd254))) begin
        tmp_V_255_fu_2278 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd255))) begin
        tmp_V_256_fu_2282 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd256))) begin
        tmp_V_257_fu_2286 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd257))) begin
        tmp_V_258_fu_2290 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd258))) begin
        tmp_V_259_fu_2294 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd24))) begin
        tmp_V_25_fu_1358 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd259))) begin
        tmp_V_260_fu_2298 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd260))) begin
        tmp_V_261_fu_2302 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd261))) begin
        tmp_V_262_fu_2306 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd262))) begin
        tmp_V_263_fu_2310 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd263))) begin
        tmp_V_264_fu_2314 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd264))) begin
        tmp_V_265_fu_2318 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd265))) begin
        tmp_V_266_fu_2322 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd266))) begin
        tmp_V_267_fu_2326 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd267))) begin
        tmp_V_268_fu_2330 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd268))) begin
        tmp_V_269_fu_2334 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd25))) begin
        tmp_V_26_fu_1362 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd269))) begin
        tmp_V_270_fu_2338 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd270))) begin
        tmp_V_271_fu_2342 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd271))) begin
        tmp_V_272_fu_2346 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd272))) begin
        tmp_V_273_fu_2350 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd273))) begin
        tmp_V_274_fu_2354 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd274))) begin
        tmp_V_275_fu_2358 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd275))) begin
        tmp_V_276_fu_2362 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd276))) begin
        tmp_V_277_fu_2366 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd277))) begin
        tmp_V_278_fu_2370 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd278))) begin
        tmp_V_279_fu_2374 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd26))) begin
        tmp_V_27_fu_1366 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd279))) begin
        tmp_V_280_fu_2378 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd280))) begin
        tmp_V_281_fu_2382 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd281))) begin
        tmp_V_282_fu_2386 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd282))) begin
        tmp_V_283_fu_2390 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd283))) begin
        tmp_V_284_fu_2394 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd284))) begin
        tmp_V_285_fu_2398 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd285))) begin
        tmp_V_286_fu_2402 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd286))) begin
        tmp_V_287_fu_2406 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd287))) begin
        tmp_V_288_fu_2410 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd288))) begin
        tmp_V_289_fu_2414 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd27))) begin
        tmp_V_28_fu_1370 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd289))) begin
        tmp_V_290_fu_2418 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd290))) begin
        tmp_V_291_fu_2422 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd291))) begin
        tmp_V_292_fu_2426 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd292))) begin
        tmp_V_293_fu_2430 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd293))) begin
        tmp_V_294_fu_2434 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd294))) begin
        tmp_V_295_fu_2438 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd295))) begin
        tmp_V_296_fu_2442 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd296))) begin
        tmp_V_297_fu_2446 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd297))) begin
        tmp_V_298_fu_2450 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd298))) begin
        tmp_V_299_fu_2454 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd28))) begin
        tmp_V_29_fu_1374 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd2))) begin
        tmp_V_2_fu_1270 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd299))) begin
        tmp_V_300_fu_2458 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd300))) begin
        tmp_V_301_fu_2462 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd301))) begin
        tmp_V_302_fu_2466 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd302))) begin
        tmp_V_303_fu_2470 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd303))) begin
        tmp_V_304_fu_2474 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd304))) begin
        tmp_V_305_fu_2478 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd305))) begin
        tmp_V_306_fu_2482 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd306))) begin
        tmp_V_307_fu_2486 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd307))) begin
        tmp_V_308_fu_2490 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd308))) begin
        tmp_V_309_fu_2494 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd29))) begin
        tmp_V_30_fu_1378 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd309))) begin
        tmp_V_310_fu_2498 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd310))) begin
        tmp_V_311_fu_2502 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd311))) begin
        tmp_V_312_fu_2506 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd312))) begin
        tmp_V_313_fu_2510 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd313))) begin
        tmp_V_314_fu_2514 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd314))) begin
        tmp_V_315_fu_2518 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd315))) begin
        tmp_V_316_fu_2522 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd316))) begin
        tmp_V_317_fu_2526 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd317))) begin
        tmp_V_318_fu_2530 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd318))) begin
        tmp_V_319_fu_2534 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd30))) begin
        tmp_V_31_fu_1382 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd319))) begin
        tmp_V_320_fu_2538 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd320))) begin
        tmp_V_321_fu_2542 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd321))) begin
        tmp_V_322_fu_2546 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd322))) begin
        tmp_V_323_fu_2550 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd323))) begin
        tmp_V_324_fu_2554 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd324))) begin
        tmp_V_325_fu_2558 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd325))) begin
        tmp_V_326_fu_2562 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd326))) begin
        tmp_V_327_fu_2566 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd327))) begin
        tmp_V_328_fu_2570 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd328))) begin
        tmp_V_329_fu_2574 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd31))) begin
        tmp_V_32_fu_1386 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd329))) begin
        tmp_V_330_fu_2578 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd330))) begin
        tmp_V_331_fu_2582 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd331))) begin
        tmp_V_332_fu_2586 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd332))) begin
        tmp_V_333_fu_2590 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd333))) begin
        tmp_V_334_fu_2594 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd334))) begin
        tmp_V_335_fu_2598 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd335))) begin
        tmp_V_336_fu_2602 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd336))) begin
        tmp_V_337_fu_2606 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd337))) begin
        tmp_V_338_fu_2610 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd338))) begin
        tmp_V_339_fu_2614 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd32))) begin
        tmp_V_33_fu_1390 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd339))) begin
        tmp_V_340_fu_2618 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd340))) begin
        tmp_V_341_fu_2622 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd341))) begin
        tmp_V_342_fu_2626 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd342))) begin
        tmp_V_343_fu_2630 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd343))) begin
        tmp_V_344_fu_2634 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd344))) begin
        tmp_V_345_fu_2638 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd345))) begin
        tmp_V_346_fu_2642 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd346))) begin
        tmp_V_347_fu_2646 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd347))) begin
        tmp_V_348_fu_2650 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd348))) begin
        tmp_V_349_fu_2654 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd33))) begin
        tmp_V_34_fu_1394 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd349))) begin
        tmp_V_350_fu_2658 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd350))) begin
        tmp_V_351_fu_2662 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd351))) begin
        tmp_V_352_fu_2666 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd352))) begin
        tmp_V_353_fu_2670 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd353))) begin
        tmp_V_354_fu_2674 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd354))) begin
        tmp_V_355_fu_2678 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd355))) begin
        tmp_V_356_fu_2682 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd356))) begin
        tmp_V_357_fu_2686 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd357))) begin
        tmp_V_358_fu_2690 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd358))) begin
        tmp_V_359_fu_2694 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd34))) begin
        tmp_V_35_fu_1398 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd359))) begin
        tmp_V_360_fu_2698 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd360))) begin
        tmp_V_361_fu_2702 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd361))) begin
        tmp_V_362_fu_2706 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd362))) begin
        tmp_V_363_fu_2710 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd363))) begin
        tmp_V_364_fu_2714 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd364))) begin
        tmp_V_365_fu_2718 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd365))) begin
        tmp_V_366_fu_2722 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd366))) begin
        tmp_V_367_fu_2726 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd367))) begin
        tmp_V_368_fu_2730 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd368))) begin
        tmp_V_369_fu_2734 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd35))) begin
        tmp_V_36_fu_1402 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd369))) begin
        tmp_V_370_fu_2738 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd370))) begin
        tmp_V_371_fu_2742 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd371))) begin
        tmp_V_372_fu_2746 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd372))) begin
        tmp_V_373_fu_2750 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd373))) begin
        tmp_V_374_fu_2754 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd374))) begin
        tmp_V_375_fu_2758 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd375))) begin
        tmp_V_376_fu_2762 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd376))) begin
        tmp_V_377_fu_2766 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd377))) begin
        tmp_V_378_fu_2770 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd378))) begin
        tmp_V_379_fu_2774 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd36))) begin
        tmp_V_37_fu_1406 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd379))) begin
        tmp_V_380_fu_2778 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd380))) begin
        tmp_V_381_fu_2782 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd381))) begin
        tmp_V_382_fu_2786 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd382))) begin
        tmp_V_383_fu_2790 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd383))) begin
        tmp_V_384_fu_2794 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd384))) begin
        tmp_V_385_fu_2798 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd385))) begin
        tmp_V_386_fu_2802 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd386))) begin
        tmp_V_387_fu_2806 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd387))) begin
        tmp_V_388_fu_2810 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd388))) begin
        tmp_V_389_fu_2814 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd37))) begin
        tmp_V_38_fu_1410 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd389))) begin
        tmp_V_390_fu_2818 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd390))) begin
        tmp_V_391_fu_2822 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd391))) begin
        tmp_V_392_fu_2826 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd392))) begin
        tmp_V_393_fu_2830 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd393))) begin
        tmp_V_394_fu_2834 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd394))) begin
        tmp_V_395_fu_2838 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd395))) begin
        tmp_V_396_fu_2842 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd396))) begin
        tmp_V_397_fu_2846 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd397))) begin
        tmp_V_398_fu_2850 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd398))) begin
        tmp_V_399_fu_2854 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd38))) begin
        tmp_V_39_fu_1414 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd399))) begin
        tmp_V_400_fu_2858 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd400))) begin
        tmp_V_401_fu_2862 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd401))) begin
        tmp_V_402_fu_2866 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd402))) begin
        tmp_V_403_fu_2870 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd403))) begin
        tmp_V_404_fu_2874 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd404))) begin
        tmp_V_405_fu_2878 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd405))) begin
        tmp_V_406_fu_2882 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd406))) begin
        tmp_V_407_fu_2886 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd407))) begin
        tmp_V_408_fu_2890 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd408))) begin
        tmp_V_409_fu_2894 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd39))) begin
        tmp_V_40_fu_1418 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd409))) begin
        tmp_V_410_fu_2898 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd410))) begin
        tmp_V_411_fu_2902 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd411))) begin
        tmp_V_412_fu_2906 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd412))) begin
        tmp_V_413_fu_2910 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd413))) begin
        tmp_V_414_fu_2914 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd414))) begin
        tmp_V_415_fu_2918 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd415))) begin
        tmp_V_416_fu_2922 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd416))) begin
        tmp_V_417_fu_2926 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd417))) begin
        tmp_V_418_fu_2930 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd418))) begin
        tmp_V_419_fu_2934 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd40))) begin
        tmp_V_41_fu_1422 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd419))) begin
        tmp_V_420_fu_2938 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd420))) begin
        tmp_V_421_fu_2942 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd421))) begin
        tmp_V_422_fu_2946 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd422))) begin
        tmp_V_423_fu_2950 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd423))) begin
        tmp_V_424_fu_2954 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd424))) begin
        tmp_V_425_fu_2958 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd425))) begin
        tmp_V_426_fu_2962 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd426))) begin
        tmp_V_427_fu_2966 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd427))) begin
        tmp_V_428_fu_2970 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd428))) begin
        tmp_V_429_fu_2974 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd41))) begin
        tmp_V_42_fu_1426 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd429))) begin
        tmp_V_430_fu_2978 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd430))) begin
        tmp_V_431_fu_2982 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd431))) begin
        tmp_V_432_fu_2986 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd432))) begin
        tmp_V_433_fu_2990 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd433))) begin
        tmp_V_434_fu_2994 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd434))) begin
        tmp_V_435_fu_2998 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd435))) begin
        tmp_V_436_fu_3002 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd436))) begin
        tmp_V_437_fu_3006 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd437))) begin
        tmp_V_438_fu_3010 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd438))) begin
        tmp_V_439_fu_3014 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd42))) begin
        tmp_V_43_fu_1430 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd439))) begin
        tmp_V_440_fu_3018 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd440))) begin
        tmp_V_441_fu_3022 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd441))) begin
        tmp_V_442_fu_3026 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd442))) begin
        tmp_V_443_fu_3030 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd443))) begin
        tmp_V_444_fu_3034 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd444))) begin
        tmp_V_445_fu_3038 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd445))) begin
        tmp_V_446_fu_3042 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd446))) begin
        tmp_V_447_fu_3046 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd447))) begin
        tmp_V_448_fu_3050 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd448))) begin
        tmp_V_449_fu_3054 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd43))) begin
        tmp_V_44_fu_1434 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd449))) begin
        tmp_V_450_fu_3058 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd450))) begin
        tmp_V_451_fu_3062 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd451))) begin
        tmp_V_452_fu_3066 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd452))) begin
        tmp_V_453_fu_3070 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd453))) begin
        tmp_V_454_fu_3074 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd454))) begin
        tmp_V_455_fu_3078 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd455))) begin
        tmp_V_456_fu_3082 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd456))) begin
        tmp_V_457_fu_3086 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd457))) begin
        tmp_V_458_fu_3090 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd458))) begin
        tmp_V_459_fu_3094 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd44))) begin
        tmp_V_45_fu_1438 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd459))) begin
        tmp_V_460_fu_3098 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd460))) begin
        tmp_V_461_fu_3102 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd461))) begin
        tmp_V_462_fu_3106 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd462))) begin
        tmp_V_463_fu_3110 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd463))) begin
        tmp_V_464_fu_3114 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd464))) begin
        tmp_V_465_fu_3118 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd465))) begin
        tmp_V_466_fu_3122 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd466))) begin
        tmp_V_467_fu_3126 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd467))) begin
        tmp_V_468_fu_3130 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd468))) begin
        tmp_V_469_fu_3134 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd45))) begin
        tmp_V_46_fu_1442 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd469))) begin
        tmp_V_470_fu_3138 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd470))) begin
        tmp_V_471_fu_3142 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd471))) begin
        tmp_V_472_fu_3146 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd472))) begin
        tmp_V_473_fu_3150 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd473))) begin
        tmp_V_474_fu_3154 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd474))) begin
        tmp_V_475_fu_3158 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd475))) begin
        tmp_V_476_fu_3162 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd476))) begin
        tmp_V_477_fu_3166 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd477))) begin
        tmp_V_478_fu_3170 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd478))) begin
        tmp_V_479_fu_3174 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd46))) begin
        tmp_V_47_fu_1446 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd479))) begin
        tmp_V_480_fu_3178 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd480))) begin
        tmp_V_481_fu_3182 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd481))) begin
        tmp_V_482_fu_3186 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd482))) begin
        tmp_V_483_fu_3190 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd483))) begin
        tmp_V_484_fu_3194 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd484))) begin
        tmp_V_485_fu_3198 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd485))) begin
        tmp_V_486_fu_3202 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd486))) begin
        tmp_V_487_fu_3206 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd487))) begin
        tmp_V_488_fu_3210 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd488))) begin
        tmp_V_489_fu_3214 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd47))) begin
        tmp_V_48_fu_1450 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd489))) begin
        tmp_V_490_fu_3218 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd490))) begin
        tmp_V_491_fu_3222 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd491))) begin
        tmp_V_492_fu_3226 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd492))) begin
        tmp_V_493_fu_3230 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd493))) begin
        tmp_V_494_fu_3234 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd494))) begin
        tmp_V_495_fu_3238 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd495))) begin
        tmp_V_496_fu_3242 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd496))) begin
        tmp_V_497_fu_3246 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd497))) begin
        tmp_V_498_fu_3250 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd498))) begin
        tmp_V_499_fu_3254 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd48))) begin
        tmp_V_49_fu_1454 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd3))) begin
        tmp_V_4_fu_1274 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd499))) begin
        tmp_V_500_fu_3258 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd500))) begin
        tmp_V_501_fu_3262 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd501))) begin
        tmp_V_502_fu_3266 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd502))) begin
        tmp_V_503_fu_3270 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd503))) begin
        tmp_V_504_fu_3274 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd504))) begin
        tmp_V_505_fu_3278 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd505))) begin
        tmp_V_506_fu_3282 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd506))) begin
        tmp_V_507_fu_3286 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd507))) begin
        tmp_V_508_fu_3290 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd508))) begin
        tmp_V_509_fu_3294 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd49))) begin
        tmp_V_50_fu_1458 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd509))) begin
        tmp_V_510_fu_3298 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd510))) begin
        tmp_V_511_fu_3302 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd511))) begin
        tmp_V_512_fu_3306 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd512))) begin
        tmp_V_513_fu_3310 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd513))) begin
        tmp_V_514_fu_3314 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd514))) begin
        tmp_V_515_fu_3318 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd515))) begin
        tmp_V_516_fu_3322 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd516))) begin
        tmp_V_517_fu_3326 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd517))) begin
        tmp_V_518_fu_3330 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd518))) begin
        tmp_V_519_fu_3334 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd50))) begin
        tmp_V_51_fu_1462 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd519))) begin
        tmp_V_520_fu_3338 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd520))) begin
        tmp_V_521_fu_3342 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd521))) begin
        tmp_V_522_fu_3346 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd522))) begin
        tmp_V_523_fu_3350 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd523))) begin
        tmp_V_524_fu_3354 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd524))) begin
        tmp_V_525_fu_3358 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd525))) begin
        tmp_V_526_fu_3362 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd526))) begin
        tmp_V_527_fu_3366 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd527))) begin
        tmp_V_528_fu_3370 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd528))) begin
        tmp_V_529_fu_3374 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd51))) begin
        tmp_V_52_fu_1466 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd529))) begin
        tmp_V_530_fu_3378 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd530))) begin
        tmp_V_531_fu_3382 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd531))) begin
        tmp_V_532_fu_3386 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd532))) begin
        tmp_V_533_fu_3390 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd533))) begin
        tmp_V_534_fu_3394 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd534))) begin
        tmp_V_535_fu_3398 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd535))) begin
        tmp_V_536_fu_3402 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd536))) begin
        tmp_V_537_fu_3406 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd537))) begin
        tmp_V_538_fu_3410 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd538))) begin
        tmp_V_539_fu_3414 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd52))) begin
        tmp_V_53_fu_1470 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd539))) begin
        tmp_V_540_fu_3418 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd540))) begin
        tmp_V_541_fu_3422 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd541))) begin
        tmp_V_542_fu_3426 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd542))) begin
        tmp_V_543_fu_3430 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd543))) begin
        tmp_V_544_fu_3434 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd544))) begin
        tmp_V_545_fu_3438 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd545))) begin
        tmp_V_546_fu_3442 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd546))) begin
        tmp_V_547_fu_3446 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd547))) begin
        tmp_V_548_fu_3450 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd548))) begin
        tmp_V_549_fu_3454 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd53))) begin
        tmp_V_54_fu_1474 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd549))) begin
        tmp_V_550_fu_3458 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd550))) begin
        tmp_V_551_fu_3462 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd551))) begin
        tmp_V_552_fu_3466 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd552))) begin
        tmp_V_553_fu_3470 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd553))) begin
        tmp_V_554_fu_3474 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd554))) begin
        tmp_V_555_fu_3478 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd555))) begin
        tmp_V_556_fu_3482 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd556))) begin
        tmp_V_557_fu_3486 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd557))) begin
        tmp_V_558_fu_3490 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd558))) begin
        tmp_V_559_fu_3494 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd54))) begin
        tmp_V_55_fu_1478 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd559))) begin
        tmp_V_560_fu_3498 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd560))) begin
        tmp_V_561_fu_3502 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd561))) begin
        tmp_V_562_fu_3506 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd562))) begin
        tmp_V_563_fu_3510 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd563))) begin
        tmp_V_564_fu_3514 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd564))) begin
        tmp_V_565_fu_3518 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd565))) begin
        tmp_V_566_fu_3522 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd566))) begin
        tmp_V_567_fu_3526 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd567))) begin
        tmp_V_568_fu_3530 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd568))) begin
        tmp_V_569_fu_3534 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd55))) begin
        tmp_V_56_fu_1482 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd569))) begin
        tmp_V_570_fu_3538 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd570))) begin
        tmp_V_571_fu_3542 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd571))) begin
        tmp_V_572_fu_3546 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd572))) begin
        tmp_V_573_fu_3550 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd573))) begin
        tmp_V_574_fu_3554 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd574))) begin
        tmp_V_575_fu_3558 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if ((~(trunc_ln321_fu_7683_p1 == 10'd214) & ~(trunc_ln321_fu_7683_p1 == 10'd213) & ~(trunc_ln321_fu_7683_p1 == 10'd212) & ~(trunc_ln321_fu_7683_p1 == 10'd211) & ~(trunc_ln321_fu_7683_p1 == 10'd210) & ~(trunc_ln321_fu_7683_p1 == 10'd209) & ~(trunc_ln321_fu_7683_p1 == 10'd208) & ~(trunc_ln321_fu_7683_p1 == 10'd207) & ~(trunc_ln321_fu_7683_p1 == 10'd206) & ~(trunc_ln321_fu_7683_p1 == 10'd205) & ~(trunc_ln321_fu_7683_p1 == 10'd204) & ~(trunc_ln321_fu_7683_p1 == 10'd203) & ~(trunc_ln321_fu_7683_p1 == 10'd202) & ~(trunc_ln321_fu_7683_p1 == 10'd201) & ~(trunc_ln321_fu_7683_p1 == 10'd200) & ~(trunc_ln321_fu_7683_p1 == 10'd199) & ~(trunc_ln321_fu_7683_p1 == 10'd198) & ~(trunc_ln321_fu_7683_p1 == 10'd197) & ~(trunc_ln321_fu_7683_p1 == 10'd196) & ~(trunc_ln321_fu_7683_p1 == 10'd195) & ~(trunc_ln321_fu_7683_p1 == 10'd194) & ~(trunc_ln321_fu_7683_p1 == 10'd193) & ~(trunc_ln321_fu_7683_p1 == 10'd192) & ~(trunc_ln321_fu_7683_p1 == 10'd191) & ~(trunc_ln321_fu_7683_p1 == 10'd190) & ~(trunc_ln321_fu_7683_p1 == 10'd189) & ~(trunc_ln321_fu_7683_p1 == 10'd188) & ~(trunc_ln321_fu_7683_p1 == 10'd187) & ~(trunc_ln321_fu_7683_p1 == 10'd186) & ~(trunc_ln321_fu_7683_p1 == 10'd185) & ~(trunc_ln321_fu_7683_p1 == 10'd184) & ~(trunc_ln321_fu_7683_p1 == 10'd183) & ~(trunc_ln321_fu_7683_p1 == 10'd182) & ~(trunc_ln321_fu_7683_p1 == 10'd181) & ~(trunc_ln321_fu_7683_p1 == 10'd180) & ~(trunc_ln321_fu_7683_p1 == 10'd179) & ~(trunc_ln321_fu_7683_p1 == 10'd178) & ~(trunc_ln321_fu_7683_p1 == 10'd177) & ~(trunc_ln321_fu_7683_p1 == 10'd176) & ~(trunc_ln321_fu_7683_p1 == 10'd175) & ~(trunc_ln321_fu_7683_p1 == 10'd174) & ~(trunc_ln321_fu_7683_p1 == 10'd173) & ~(trunc_ln321_fu_7683_p1 == 10'd172) & ~(trunc_ln321_fu_7683_p1 == 10'd171) & ~(trunc_ln321_fu_7683_p1 == 10'd170) & ~(trunc_ln321_fu_7683_p1 == 10'd169) & ~(trunc_ln321_fu_7683_p1 == 10'd168) & ~(trunc_ln321_fu_7683_p1 == 10'd167) & ~(trunc_ln321_fu_7683_p1 == 10'd166) & ~(trunc_ln321_fu_7683_p1 == 10'd165) & ~(trunc_ln321_fu_7683_p1 == 10'd164) & ~(trunc_ln321_fu_7683_p1 == 10'd163) & ~(trunc_ln321_fu_7683_p1 == 10'd162) & ~(trunc_ln321_fu_7683_p1 == 10'd161) & ~(trunc_ln321_fu_7683_p1 == 10'd160) & ~(trunc_ln321_fu_7683_p1 == 10'd159) & ~(trunc_ln321_fu_7683_p1 == 10'd158) & ~(trunc_ln321_fu_7683_p1 == 10'd157) & ~(trunc_ln321_fu_7683_p1 == 10'd156) & ~(trunc_ln321_fu_7683_p1 == 10'd155) & ~(trunc_ln321_fu_7683_p1 == 10'd154) & ~(trunc_ln321_fu_7683_p1 == 10'd153) & ~(trunc_ln321_fu_7683_p1 == 10'd152) & ~(trunc_ln321_fu_7683_p1 == 10'd151) & ~(trunc_ln321_fu_7683_p1 == 10'd150) & ~(trunc_ln321_fu_7683_p1 == 10'd149) & ~(trunc_ln321_fu_7683_p1 == 10'd148) & ~(trunc_ln321_fu_7683_p1 == 10'd147) & ~(trunc_ln321_fu_7683_p1 == 10'd146) & ~(trunc_ln321_fu_7683_p1 == 10'd145) & ~(trunc_ln321_fu_7683_p1 == 10'd144) & ~(trunc_ln321_fu_7683_p1 == 10'd143) & ~(trunc_ln321_fu_7683_p1 == 10'd142) & ~(trunc_ln321_fu_7683_p1 == 10'd141) & ~(trunc_ln321_fu_7683_p1 == 10'd140) & ~(trunc_ln321_fu_7683_p1 == 10'd139) & ~(trunc_ln321_fu_7683_p1 == 10'd138) & ~(trunc_ln321_fu_7683_p1 == 10'd137) & ~(trunc_ln321_fu_7683_p1 == 10'd136) & ~(trunc_ln321_fu_7683_p1 == 10'd135) & ~(trunc_ln321_fu_7683_p1 == 10'd134) & ~(trunc_ln321_fu_7683_p1 == 10'd133) & ~(trunc_ln321_fu_7683_p1 == 10'd132) & ~(trunc_ln321_fu_7683_p1 == 10'd131) & ~(trunc_ln321_fu_7683_p1 == 10'd130) & ~(trunc_ln321_fu_7683_p1 == 10'd129) & ~(trunc_ln321_fu_7683_p1 == 10'd128) & ~(trunc_ln321_fu_7683_p1 == 10'd127) & ~(trunc_ln321_fu_7683_p1 == 10'd126) & ~(trunc_ln321_fu_7683_p1 == 10'd125) & ~(trunc_ln321_fu_7683_p1 == 10'd124) & ~(trunc_ln321_fu_7683_p1 == 10'd123) & ~(trunc_ln321_fu_7683_p1 == 10'd122) & ~(trunc_ln321_fu_7683_p1 == 10'd121) & ~(trunc_ln321_fu_7683_p1 == 10'd120) & ~(trunc_ln321_fu_7683_p1 == 10'd119) & ~(trunc_ln321_fu_7683_p1 == 10'd118) & ~(trunc_ln321_fu_7683_p1 == 10'd117) & ~(trunc_ln321_fu_7683_p1 == 10'd116) & ~(trunc_ln321_fu_7683_p1 == 10'd115) & ~(trunc_ln321_fu_7683_p1 == 10'd114) & ~(trunc_ln321_fu_7683_p1 == 10'd113) & ~(trunc_ln321_fu_7683_p1 == 10'd112) & ~(trunc_ln321_fu_7683_p1 == 10'd111) & ~(trunc_ln321_fu_7683_p1 == 10'd110) & ~(trunc_ln321_fu_7683_p1 == 10'd109) & ~(trunc_ln321_fu_7683_p1 == 10'd108) & ~(trunc_ln321_fu_7683_p1 == 10'd107) & ~(trunc_ln321_fu_7683_p1 == 10'd106) & ~(trunc_ln321_fu_7683_p1 == 10'd105) & ~(trunc_ln321_fu_7683_p1 == 10'd104) & ~(trunc_ln321_fu_7683_p1 == 10'd103) & ~(trunc_ln321_fu_7683_p1 == 10'd102) & ~(trunc_ln321_fu_7683_p1 == 10'd101) & ~(trunc_ln321_fu_7683_p1 == 10'd100) & ~(trunc_ln321_fu_7683_p1 == 10'd99) & ~(trunc_ln321_fu_7683_p1 == 10'd98) & ~(trunc_ln321_fu_7683_p1 == 10'd97) & ~(trunc_ln321_fu_7683_p1 == 10'd96) & ~(trunc_ln321_fu_7683_p1 == 10'd95) & ~(trunc_ln321_fu_7683_p1 == 10'd94) & ~(trunc_ln321_fu_7683_p1 == 10'd93) & ~(trunc_ln321_fu_7683_p1 == 10'd92) & ~(trunc_ln321_fu_7683_p1 == 10'd91) & ~(trunc_ln321_fu_7683_p1 == 10'd90) & ~(trunc_ln321_fu_7683_p1 == 10'd89) & ~(trunc_ln321_fu_7683_p1 == 10'd88) & ~(trunc_ln321_fu_7683_p1 == 10'd87) & ~(trunc_ln321_fu_7683_p1 == 10'd86) & ~(trunc_ln321_fu_7683_p1 == 10'd85) & ~(trunc_ln321_fu_7683_p1 == 10'd84) & ~(trunc_ln321_fu_7683_p1 == 10'd83) & ~(trunc_ln321_fu_7683_p1 == 10'd82) & ~(trunc_ln321_fu_7683_p1 == 10'd81) & ~(trunc_ln321_fu_7683_p1 == 10'd80) & ~(trunc_ln321_fu_7683_p1 == 10'd79) & ~(trunc_ln321_fu_7683_p1 == 10'd78) & ~(trunc_ln321_fu_7683_p1 == 10'd77) & ~(trunc_ln321_fu_7683_p1 == 10'd76) & ~(trunc_ln321_fu_7683_p1 == 10'd75) & ~(trunc_ln321_fu_7683_p1 == 10'd74) & ~(trunc_ln321_fu_7683_p1 == 10'd73) & ~(trunc_ln321_fu_7683_p1 == 10'd72) & ~(trunc_ln321_fu_7683_p1 == 10'd71) & ~(trunc_ln321_fu_7683_p1 == 10'd70) & ~(trunc_ln321_fu_7683_p1 == 10'd69) & ~(trunc_ln321_fu_7683_p1 == 10'd68) & ~(trunc_ln321_fu_7683_p1 == 10'd67) & ~(trunc_ln321_fu_7683_p1 == 10'd66) & ~(trunc_ln321_fu_7683_p1 == 10'd65) & ~(trunc_ln321_fu_7683_p1 == 10'd64) & ~(trunc_ln321_fu_7683_p1 == 10'd63) & ~(trunc_ln321_fu_7683_p1 == 10'd62) & ~(trunc_ln321_fu_7683_p1 == 10'd61) & ~(trunc_ln321_fu_7683_p1 == 10'd60) & ~(trunc_ln321_fu_7683_p1 == 10'd59) & ~(trunc_ln321_fu_7683_p1 == 10'd58) & ~(trunc_ln321_fu_7683_p1 == 10'd57) & ~(trunc_ln321_fu_7683_p1 == 10'd56) & ~(trunc_ln321_fu_7683_p1 == 10'd55) & ~(trunc_ln321_fu_7683_p1 == 10'd54) & ~(trunc_ln321_fu_7683_p1 == 10'd53) & ~(trunc_ln321_fu_7683_p1 == 10'd52) & ~(trunc_ln321_fu_7683_p1 == 10'd51) & ~(trunc_ln321_fu_7683_p1 == 10'd50) & ~(trunc_ln321_fu_7683_p1 == 10'd49) & ~(trunc_ln321_fu_7683_p1 == 10'd48) & ~(trunc_ln321_fu_7683_p1 == 10'd47) & ~(trunc_ln321_fu_7683_p1 == 10'd46) & ~(trunc_ln321_fu_7683_p1 == 10'd45) & ~(trunc_ln321_fu_7683_p1 == 10'd44) & ~(trunc_ln321_fu_7683_p1 == 10'd43) & ~(trunc_ln321_fu_7683_p1 == 10'd42) & ~(trunc_ln321_fu_7683_p1 == 10'd41) & ~(trunc_ln321_fu_7683_p1 == 10'd40) & ~(trunc_ln321_fu_7683_p1 == 10'd39) & ~(trunc_ln321_fu_7683_p1 == 10'd38) & ~(trunc_ln321_fu_7683_p1 == 10'd37) & ~(trunc_ln321_fu_7683_p1 == 10'd36) & ~(trunc_ln321_fu_7683_p1 == 10'd35) & ~(trunc_ln321_fu_7683_p1 == 10'd34) & ~(trunc_ln321_fu_7683_p1 == 10'd33) & ~(trunc_ln321_fu_7683_p1 == 10'd32) & ~(trunc_ln321_fu_7683_p1 == 10'd31) & ~(trunc_ln321_fu_7683_p1 == 10'd30) & ~(trunc_ln321_fu_7683_p1 == 10'd29) & ~(trunc_ln321_fu_7683_p1 == 10'd28) & ~(trunc_ln321_fu_7683_p1 == 10'd27) & ~(trunc_ln321_fu_7683_p1 == 10'd26) & ~(trunc_ln321_fu_7683_p1 == 10'd574) & ~(trunc_ln321_fu_7683_p1 == 10'd573) & ~(trunc_ln321_fu_7683_p1 == 10'd572) & ~(trunc_ln321_fu_7683_p1 == 10'd25) & ~(trunc_ln321_fu_7683_p1 == 10'd571) & ~(trunc_ln321_fu_7683_p1 == 10'd570) & ~(trunc_ln321_fu_7683_p1 == 10'd569) & ~(trunc_ln321_fu_7683_p1 == 10'd568) & ~(trunc_ln321_fu_7683_p1 == 10'd567) & ~(trunc_ln321_fu_7683_p1 == 10'd566) & ~(trunc_ln321_fu_7683_p1 == 10'd565) & ~(trunc_ln321_fu_7683_p1 == 10'd564) & ~(trunc_ln321_fu_7683_p1 == 10'd563) & ~(trunc_ln321_fu_7683_p1 == 10'd562) & ~(trunc_ln321_fu_7683_p1 == 10'd24) & ~(trunc_ln321_fu_7683_p1 == 10'd561) & ~(trunc_ln321_fu_7683_p1 == 10'd560) & ~(trunc_ln321_fu_7683_p1 == 10'd559) & ~(trunc_ln321_fu_7683_p1 == 10'd558) & ~(trunc_ln321_fu_7683_p1 == 10'd557) & ~(trunc_ln321_fu_7683_p1 == 10'd556) & ~(trunc_ln321_fu_7683_p1 == 10'd555) & ~(trunc_ln321_fu_7683_p1 == 10'd554) & ~(trunc_ln321_fu_7683_p1 == 10'd553) & ~(trunc_ln321_fu_7683_p1 == 10'd552) & ~(trunc_ln321_fu_7683_p1 == 10'd23) & ~(trunc_ln321_fu_7683_p1 == 10'd551) & ~(trunc_ln321_fu_7683_p1 == 10'd550) & ~(trunc_ln321_fu_7683_p1 == 10'd549) & ~(trunc_ln321_fu_7683_p1 == 10'd548) & ~(trunc_ln321_fu_7683_p1 == 10'd547) & ~(trunc_ln321_fu_7683_p1 == 10'd546) & ~(trunc_ln321_fu_7683_p1 == 10'd545) & ~(trunc_ln321_fu_7683_p1 == 10'd544) & ~(trunc_ln321_fu_7683_p1 == 10'd543) & ~(trunc_ln321_fu_7683_p1 == 10'd542) & ~(trunc_ln321_fu_7683_p1 == 10'd22) & ~(trunc_ln321_fu_7683_p1 == 10'd541) & ~(trunc_ln321_fu_7683_p1 == 10'd540) & ~(trunc_ln321_fu_7683_p1 == 10'd539) & ~(trunc_ln321_fu_7683_p1 == 10'd538) & ~(trunc_ln321_fu_7683_p1 == 10'd537) & ~(trunc_ln321_fu_7683_p1 == 10'd536) & ~(trunc_ln321_fu_7683_p1 == 10'd535) & ~(trunc_ln321_fu_7683_p1 == 10'd534) & ~(trunc_ln321_fu_7683_p1 == 10'd533) & ~(trunc_ln321_fu_7683_p1 == 10'd532) & ~(trunc_ln321_fu_7683_p1 == 10'd21) & ~(trunc_ln321_fu_7683_p1 == 10'd531) & ~(trunc_ln321_fu_7683_p1 == 10'd530) & ~(trunc_ln321_fu_7683_p1 == 10'd529) & ~(trunc_ln321_fu_7683_p1 == 10'd528) & ~(trunc_ln321_fu_7683_p1 == 10'd527) & ~(trunc_ln321_fu_7683_p1 == 10'd526) & ~(trunc_ln321_fu_7683_p1 == 10'd525) & ~(trunc_ln321_fu_7683_p1 == 10'd524) & ~(trunc_ln321_fu_7683_p1 == 10'd523) & ~(trunc_ln321_fu_7683_p1 == 10'd522) & ~(trunc_ln321_fu_7683_p1 == 10'd20) & ~(trunc_ln321_fu_7683_p1 == 10'd521) & ~(trunc_ln321_fu_7683_p1 == 10'd520) & ~(trunc_ln321_fu_7683_p1 == 10'd519) & ~(trunc_ln321_fu_7683_p1 == 10'd518) & ~(trunc_ln321_fu_7683_p1 == 10'd517) & ~(trunc_ln321_fu_7683_p1 == 10'd516) & ~(trunc_ln321_fu_7683_p1 == 10'd515) & ~(trunc_ln321_fu_7683_p1 == 10'd514) & ~(trunc_ln321_fu_7683_p1 == 10'd513) & ~(trunc_ln321_fu_7683_p1 == 10'd512) & ~(trunc_ln321_fu_7683_p1 == 10'd19) & ~(trunc_ln321_fu_7683_p1 == 10'd511) & ~(trunc_ln321_fu_7683_p1 == 10'd510) & ~(trunc_ln321_fu_7683_p1 == 10'd509) & ~(trunc_ln321_fu_7683_p1 == 10'd508) & ~(trunc_ln321_fu_7683_p1 == 10'd507) & ~(trunc_ln321_fu_7683_p1 == 10'd506) & ~(trunc_ln321_fu_7683_p1 == 10'd505) & ~(trunc_ln321_fu_7683_p1 == 10'd504) & ~(trunc_ln321_fu_7683_p1 == 10'd503) & ~(trunc_ln321_fu_7683_p1 == 10'd502) & ~(trunc_ln321_fu_7683_p1 == 10'd18) & ~(trunc_ln321_fu_7683_p1 == 10'd501) & ~(trunc_ln321_fu_7683_p1 == 10'd500) & ~(trunc_ln321_fu_7683_p1 == 10'd499) & ~(trunc_ln321_fu_7683_p1 == 10'd498) & ~(trunc_ln321_fu_7683_p1 == 10'd497) & ~(trunc_ln321_fu_7683_p1 == 10'd496) & ~(trunc_ln321_fu_7683_p1 == 10'd495) & ~(trunc_ln321_fu_7683_p1 == 10'd494) & ~(trunc_ln321_fu_7683_p1 == 10'd493) & ~(trunc_ln321_fu_7683_p1 == 10'd492) & ~(trunc_ln321_fu_7683_p1 == 10'd17) & ~(trunc_ln321_fu_7683_p1 == 10'd491) & ~(trunc_ln321_fu_7683_p1 == 10'd490) & ~(trunc_ln321_fu_7683_p1 == 10'd489) & ~(trunc_ln321_fu_7683_p1 == 10'd488) & ~(trunc_ln321_fu_7683_p1 == 10'd487) & ~(trunc_ln321_fu_7683_p1 == 10'd486) & ~(trunc_ln321_fu_7683_p1 == 10'd485) & ~(trunc_ln321_fu_7683_p1 == 10'd484) & ~(trunc_ln321_fu_7683_p1 == 10'd483) & ~(trunc_ln321_fu_7683_p1 == 10'd482) & ~(trunc_ln321_fu_7683_p1 == 10'd16) & ~(trunc_ln321_fu_7683_p1 == 10'd481) & ~(trunc_ln321_fu_7683_p1 == 10'd480) & ~(trunc_ln321_fu_7683_p1 == 10'd479) & ~(trunc_ln321_fu_7683_p1 == 10'd478) & ~(trunc_ln321_fu_7683_p1 == 10'd477) & ~(trunc_ln321_fu_7683_p1 == 10'd476) & ~(trunc_ln321_fu_7683_p1 == 10'd475) & ~(trunc_ln321_fu_7683_p1 == 10'd474) & ~(trunc_ln321_fu_7683_p1 == 10'd473) & ~(trunc_ln321_fu_7683_p1 == 10'd472) & ~(trunc_ln321_fu_7683_p1 == 10'd15) & ~(trunc_ln321_fu_7683_p1 == 10'd471) & ~(trunc_ln321_fu_7683_p1 == 10'd470) & ~(trunc_ln321_fu_7683_p1 == 10'd469) & ~(trunc_ln321_fu_7683_p1 == 10'd468) & ~(trunc_ln321_fu_7683_p1 == 10'd467) & ~(trunc_ln321_fu_7683_p1 == 10'd466) & ~(trunc_ln321_fu_7683_p1 == 10'd465) & ~(trunc_ln321_fu_7683_p1 == 10'd464) & ~(trunc_ln321_fu_7683_p1 == 10'd463) & ~(trunc_ln321_fu_7683_p1 == 10'd462) & ~(trunc_ln321_fu_7683_p1 == 10'd14) & ~(trunc_ln321_fu_7683_p1 == 10'd461) & ~(trunc_ln321_fu_7683_p1 == 10'd460) & ~(trunc_ln321_fu_7683_p1 == 10'd459) & ~(trunc_ln321_fu_7683_p1 == 10'd458) & ~(trunc_ln321_fu_7683_p1 == 10'd457) & ~(trunc_ln321_fu_7683_p1 == 10'd456) & ~(trunc_ln321_fu_7683_p1 == 10'd455) & ~(trunc_ln321_fu_7683_p1 == 10'd454) & ~(trunc_ln321_fu_7683_p1 == 10'd453) & ~(trunc_ln321_fu_7683_p1 == 10'd452) & ~(trunc_ln321_fu_7683_p1 == 10'd13) & ~(trunc_ln321_fu_7683_p1 == 10'd451) & ~(trunc_ln321_fu_7683_p1 == 10'd450) & ~(trunc_ln321_fu_7683_p1 == 10'd449) & ~(trunc_ln321_fu_7683_p1 == 10'd448) & ~(trunc_ln321_fu_7683_p1 == 10'd447) & ~(trunc_ln321_fu_7683_p1 == 10'd446) & ~(trunc_ln321_fu_7683_p1 == 10'd445) & ~(trunc_ln321_fu_7683_p1 == 10'd444) & ~(trunc_ln321_fu_7683_p1 == 10'd443) & ~(trunc_ln321_fu_7683_p1 == 10'd442) & ~(trunc_ln321_fu_7683_p1 == 10'd12) & ~(trunc_ln321_fu_7683_p1 == 10'd441) & ~(trunc_ln321_fu_7683_p1 == 10'd440) & ~(trunc_ln321_fu_7683_p1 == 10'd439) & ~(trunc_ln321_fu_7683_p1 == 10'd438) & ~(trunc_ln321_fu_7683_p1 == 10'd437) & ~(trunc_ln321_fu_7683_p1 == 10'd436) & ~(trunc_ln321_fu_7683_p1 == 10'd435) & ~(trunc_ln321_fu_7683_p1 == 10'd434) & ~(trunc_ln321_fu_7683_p1 == 10'd433) & ~(trunc_ln321_fu_7683_p1 == 10'd432) & ~(trunc_ln321_fu_7683_p1 == 10'd11) & ~(trunc_ln321_fu_7683_p1 == 10'd431) & ~(trunc_ln321_fu_7683_p1 == 10'd430) & ~(trunc_ln321_fu_7683_p1 == 10'd429) & ~(trunc_ln321_fu_7683_p1 == 10'd428) & ~(trunc_ln321_fu_7683_p1 == 10'd427) & ~(trunc_ln321_fu_7683_p1 == 10'd426) & ~(trunc_ln321_fu_7683_p1 == 10'd425) & ~(trunc_ln321_fu_7683_p1 == 10'd424) & ~(trunc_ln321_fu_7683_p1 == 10'd423) & ~(trunc_ln321_fu_7683_p1 == 10'd422) & ~(trunc_ln321_fu_7683_p1 == 10'd10) & ~(trunc_ln321_fu_7683_p1 == 10'd421) & ~(trunc_ln321_fu_7683_p1 == 10'd420) & ~(trunc_ln321_fu_7683_p1 == 10'd419) & ~(trunc_ln321_fu_7683_p1 == 10'd418) & ~(trunc_ln321_fu_7683_p1 == 10'd417) & ~(trunc_ln321_fu_7683_p1 == 10'd416) & ~(trunc_ln321_fu_7683_p1 == 10'd415) & ~(trunc_ln321_fu_7683_p1 == 10'd414) & ~(trunc_ln321_fu_7683_p1 == 10'd413) & ~(trunc_ln321_fu_7683_p1 == 10'd412) & ~(trunc_ln321_fu_7683_p1 == 10'd9) & ~(trunc_ln321_fu_7683_p1 == 10'd411) & ~(trunc_ln321_fu_7683_p1 == 10'd410) & ~(trunc_ln321_fu_7683_p1 == 10'd409) & ~(trunc_ln321_fu_7683_p1 == 10'd408) & ~(trunc_ln321_fu_7683_p1 == 10'd407) & ~(trunc_ln321_fu_7683_p1 == 10'd406) & ~(trunc_ln321_fu_7683_p1 == 10'd405) & ~(trunc_ln321_fu_7683_p1 == 10'd404) & ~(trunc_ln321_fu_7683_p1 == 10'd403) & ~(trunc_ln321_fu_7683_p1 == 10'd402) & ~(trunc_ln321_fu_7683_p1 == 10'd8) & ~(trunc_ln321_fu_7683_p1 == 10'd401) & ~(trunc_ln321_fu_7683_p1 == 10'd400) & ~(trunc_ln321_fu_7683_p1 == 10'd399) & ~(trunc_ln321_fu_7683_p1 == 10'd398) & ~(trunc_ln321_fu_7683_p1 == 10'd397) & ~(trunc_ln321_fu_7683_p1 == 10'd396) & ~(trunc_ln321_fu_7683_p1 == 10'd395) & ~(trunc_ln321_fu_7683_p1 == 10'd394) & ~(trunc_ln321_fu_7683_p1 == 10'd393) & ~(trunc_ln321_fu_7683_p1 == 10'd392) & ~(trunc_ln321_fu_7683_p1 == 10'd7) & ~(trunc_ln321_fu_7683_p1 == 10'd391) & ~(trunc_ln321_fu_7683_p1 == 10'd390) & ~(trunc_ln321_fu_7683_p1 == 10'd389) & ~(trunc_ln321_fu_7683_p1 == 10'd388) & ~(trunc_ln321_fu_7683_p1 == 10'd387) & ~(trunc_ln321_fu_7683_p1 == 10'd386) & ~(trunc_ln321_fu_7683_p1 == 10'd385) & ~(trunc_ln321_fu_7683_p1 == 10'd384) & ~(trunc_ln321_fu_7683_p1 == 10'd383) & ~(trunc_ln321_fu_7683_p1 == 10'd382) & ~(trunc_ln321_fu_7683_p1 == 10'd6) & ~(trunc_ln321_fu_7683_p1 == 10'd381) & ~(trunc_ln321_fu_7683_p1 == 10'd380) & ~(trunc_ln321_fu_7683_p1 == 10'd379) & ~(trunc_ln321_fu_7683_p1 == 10'd378) & ~(trunc_ln321_fu_7683_p1 == 10'd377) & ~(trunc_ln321_fu_7683_p1 == 10'd376) & ~(trunc_ln321_fu_7683_p1 == 10'd375) & ~(trunc_ln321_fu_7683_p1 == 10'd374) & ~(trunc_ln321_fu_7683_p1 == 10'd373) & ~(trunc_ln321_fu_7683_p1 == 10'd372) & ~(trunc_ln321_fu_7683_p1 == 10'd5) & ~(trunc_ln321_fu_7683_p1 == 10'd371) & ~(trunc_ln321_fu_7683_p1 == 10'd370) & ~(trunc_ln321_fu_7683_p1 == 10'd369) & ~(trunc_ln321_fu_7683_p1 == 10'd368) & ~(trunc_ln321_fu_7683_p1 == 10'd367) & ~(trunc_ln321_fu_7683_p1 == 10'd366) & ~(trunc_ln321_fu_7683_p1 == 10'd365) & ~(trunc_ln321_fu_7683_p1 == 10'd364) & ~(trunc_ln321_fu_7683_p1 == 10'd363) & ~(trunc_ln321_fu_7683_p1 == 10'd362) & ~(trunc_ln321_fu_7683_p1 == 10'd4) & ~(trunc_ln321_fu_7683_p1 == 10'd361) & ~(trunc_ln321_fu_7683_p1 == 10'd360) & ~(trunc_ln321_fu_7683_p1 == 10'd359) & ~(trunc_ln321_fu_7683_p1 == 10'd358) & ~(trunc_ln321_fu_7683_p1 == 10'd357) & ~(trunc_ln321_fu_7683_p1 == 10'd356) & ~(trunc_ln321_fu_7683_p1 == 10'd355) & ~(trunc_ln321_fu_7683_p1 == 10'd354) & ~(trunc_ln321_fu_7683_p1 == 10'd353) & ~(trunc_ln321_fu_7683_p1 == 10'd352) & ~(trunc_ln321_fu_7683_p1 == 10'd3) & ~(trunc_ln321_fu_7683_p1 == 10'd351) & ~(trunc_ln321_fu_7683_p1 == 10'd350) & ~(trunc_ln321_fu_7683_p1 == 10'd349) & ~(trunc_ln321_fu_7683_p1 == 10'd348) & ~(trunc_ln321_fu_7683_p1 == 10'd347) & ~(trunc_ln321_fu_7683_p1 == 10'd346) & ~(trunc_ln321_fu_7683_p1 == 10'd345) & ~(trunc_ln321_fu_7683_p1 == 10'd344) & ~(trunc_ln321_fu_7683_p1 == 10'd343) & ~(trunc_ln321_fu_7683_p1 == 10'd342) & ~(trunc_ln321_fu_7683_p1 == 10'd2) & ~(trunc_ln321_fu_7683_p1 == 10'd341) & ~(trunc_ln321_fu_7683_p1 == 10'd340) & ~(trunc_ln321_fu_7683_p1 == 10'd339) & ~(trunc_ln321_fu_7683_p1 == 10'd338) & ~(trunc_ln321_fu_7683_p1 == 10'd337) & ~(trunc_ln321_fu_7683_p1 == 10'd336) & ~(trunc_ln321_fu_7683_p1 == 10'd335) & ~(trunc_ln321_fu_7683_p1 == 10'd334) & ~(trunc_ln321_fu_7683_p1 == 10'd333) & ~(trunc_ln321_fu_7683_p1 == 10'd332) & ~(trunc_ln321_fu_7683_p1 == 10'd1) & ~(trunc_ln321_fu_7683_p1 == 10'd331) & ~(trunc_ln321_fu_7683_p1 == 10'd330) & ~(trunc_ln321_fu_7683_p1 == 10'd329) & ~(trunc_ln321_fu_7683_p1 == 10'd328) & ~(trunc_ln321_fu_7683_p1 == 10'd327) & ~(trunc_ln321_fu_7683_p1 == 10'd326) & ~(trunc_ln321_fu_7683_p1 == 10'd325) & ~(trunc_ln321_fu_7683_p1 == 10'd324) & ~(trunc_ln321_fu_7683_p1 == 10'd323) & ~(trunc_ln321_fu_7683_p1 == 10'd322) & ~(trunc_ln321_fu_7683_p1 == 10'd0) & ~(trunc_ln321_fu_7683_p1 == 10'd321) & ~(trunc_ln321_fu_7683_p1 == 10'd320) & ~(trunc_ln321_fu_7683_p1 == 10'd319) & ~(trunc_ln321_fu_7683_p1 == 10'd318) & ~(trunc_ln321_fu_7683_p1 == 10'd317) & ~(trunc_ln321_fu_7683_p1 == 10'd316) & ~(trunc_ln321_fu_7683_p1 == 10'd315) & ~(trunc_ln321_fu_7683_p1 == 10'd314) & ~(trunc_ln321_fu_7683_p1 == 10'd313) & ~(trunc_ln321_fu_7683_p1 == 10'd312) & ~(trunc_ln321_fu_7683_p1 == 10'd311) & ~(trunc_ln321_fu_7683_p1 == 10'd310) & ~(trunc_ln321_fu_7683_p1 == 10'd309) & ~(trunc_ln321_fu_7683_p1 == 10'd308) & ~(trunc_ln321_fu_7683_p1 == 10'd307) & ~(trunc_ln321_fu_7683_p1 == 10'd306) & ~(trunc_ln321_fu_7683_p1 == 10'd305) & ~(trunc_ln321_fu_7683_p1 == 10'd304) & ~(trunc_ln321_fu_7683_p1 == 10'd303) & ~(trunc_ln321_fu_7683_p1 == 10'd302) & ~(trunc_ln321_fu_7683_p1 == 10'd301) & ~(trunc_ln321_fu_7683_p1 == 10'd300) & ~(trunc_ln321_fu_7683_p1 == 10'd299) & ~(trunc_ln321_fu_7683_p1 == 10'd298) & ~(trunc_ln321_fu_7683_p1 == 10'd297) & ~(trunc_ln321_fu_7683_p1 == 10'd296) & ~(trunc_ln321_fu_7683_p1 == 10'd295) & ~(trunc_ln321_fu_7683_p1 == 10'd294) & ~(trunc_ln321_fu_7683_p1 == 10'd293) & ~(trunc_ln321_fu_7683_p1 == 10'd292) & ~(trunc_ln321_fu_7683_p1 == 10'd291) & ~(trunc_ln321_fu_7683_p1 == 10'd290) & ~(trunc_ln321_fu_7683_p1 == 10'd289) & ~(trunc_ln321_fu_7683_p1 == 10'd288) & ~(trunc_ln321_fu_7683_p1 == 10'd287) & ~(trunc_ln321_fu_7683_p1 == 10'd286) & ~(trunc_ln321_fu_7683_p1 == 10'd285) & ~(trunc_ln321_fu_7683_p1 == 10'd284) & ~(trunc_ln321_fu_7683_p1 == 10'd283) & ~(trunc_ln321_fu_7683_p1 == 10'd282) & ~(trunc_ln321_fu_7683_p1 == 10'd281) & ~(trunc_ln321_fu_7683_p1 == 10'd280) & ~(trunc_ln321_fu_7683_p1 == 10'd279) & ~(trunc_ln321_fu_7683_p1 == 10'd278) & ~(trunc_ln321_fu_7683_p1 == 10'd277) & ~(trunc_ln321_fu_7683_p1 == 10'd276) & ~(trunc_ln321_fu_7683_p1 == 10'd275) & ~(trunc_ln321_fu_7683_p1 == 10'd274) & ~(trunc_ln321_fu_7683_p1 == 10'd273) & ~(trunc_ln321_fu_7683_p1 == 10'd272) & ~(trunc_ln321_fu_7683_p1 == 10'd271) & ~(trunc_ln321_fu_7683_p1 == 10'd270) & ~(trunc_ln321_fu_7683_p1 == 10'd269) & ~(trunc_ln321_fu_7683_p1 == 10'd268) & ~(trunc_ln321_fu_7683_p1 == 10'd267) & ~(trunc_ln321_fu_7683_p1 == 10'd266) & ~(trunc_ln321_fu_7683_p1 == 10'd265) & ~(trunc_ln321_fu_7683_p1 == 10'd264) & ~(trunc_ln321_fu_7683_p1 == 10'd263) & ~(trunc_ln321_fu_7683_p1 == 10'd262) & ~(trunc_ln321_fu_7683_p1 == 10'd261) & ~(trunc_ln321_fu_7683_p1 == 10'd260) & ~(trunc_ln321_fu_7683_p1 == 10'd259) & ~(trunc_ln321_fu_7683_p1 == 10'd258) & ~(trunc_ln321_fu_7683_p1 == 10'd257) & ~(trunc_ln321_fu_7683_p1 == 10'd256) & ~(trunc_ln321_fu_7683_p1 == 10'd255) & ~(trunc_ln321_fu_7683_p1 == 10'd254) & ~(trunc_ln321_fu_7683_p1 == 10'd253) & ~(trunc_ln321_fu_7683_p1 == 10'd252) & ~(trunc_ln321_fu_7683_p1 == 10'd251) & ~(trunc_ln321_fu_7683_p1 == 10'd250) & ~(trunc_ln321_fu_7683_p1 == 10'd249) & ~(trunc_ln321_fu_7683_p1 == 10'd248) & ~(trunc_ln321_fu_7683_p1 == 10'd247) & ~(trunc_ln321_fu_7683_p1 == 10'd246) & ~(trunc_ln321_fu_7683_p1 == 10'd245) & ~(trunc_ln321_fu_7683_p1 == 10'd244) & ~(trunc_ln321_fu_7683_p1 == 10'd243) & ~(trunc_ln321_fu_7683_p1 == 10'd242) & ~(trunc_ln321_fu_7683_p1 == 10'd241) & ~(trunc_ln321_fu_7683_p1 == 10'd240) & ~(trunc_ln321_fu_7683_p1 == 10'd239) & ~(trunc_ln321_fu_7683_p1 == 10'd238) & ~(trunc_ln321_fu_7683_p1 == 10'd237) & ~(trunc_ln321_fu_7683_p1 == 10'd236) & ~(trunc_ln321_fu_7683_p1 == 10'd235) & ~(trunc_ln321_fu_7683_p1 == 10'd234) & ~(trunc_ln321_fu_7683_p1 == 10'd233) & ~(trunc_ln321_fu_7683_p1 == 10'd232) & ~(trunc_ln321_fu_7683_p1 == 10'd231) & ~(trunc_ln321_fu_7683_p1 == 10'd230) & ~(trunc_ln321_fu_7683_p1 == 10'd229) & ~(trunc_ln321_fu_7683_p1 == 10'd228) & ~(trunc_ln321_fu_7683_p1 == 10'd227) & ~(trunc_ln321_fu_7683_p1 == 10'd226) & ~(trunc_ln321_fu_7683_p1 == 10'd225) & ~(trunc_ln321_fu_7683_p1 == 10'd224) & ~(trunc_ln321_fu_7683_p1 == 10'd223) & ~(trunc_ln321_fu_7683_p1 == 10'd222) & ~(trunc_ln321_fu_7683_p1 == 10'd221) & ~(trunc_ln321_fu_7683_p1 == 10'd220) & ~(trunc_ln321_fu_7683_p1 == 10'd219) & ~(trunc_ln321_fu_7683_p1 == 10'd218) & ~(trunc_ln321_fu_7683_p1 == 10'd217) & ~(trunc_ln321_fu_7683_p1 == 10'd216) & ~(trunc_ln321_fu_7683_p1 == 10'd215) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_576_fu_3562 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd56))) begin
        tmp_V_57_fu_1486 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd57))) begin
        tmp_V_58_fu_1490 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd58))) begin
        tmp_V_59_fu_1494 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd4))) begin
        tmp_V_5_fu_1278 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd59))) begin
        tmp_V_60_fu_1498 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd60))) begin
        tmp_V_61_fu_1502 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd61))) begin
        tmp_V_62_fu_1506 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd62))) begin
        tmp_V_63_fu_1510 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd63))) begin
        tmp_V_64_fu_1514 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd64))) begin
        tmp_V_65_fu_1518 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd65))) begin
        tmp_V_66_fu_1522 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd66))) begin
        tmp_V_67_fu_1526 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd67))) begin
        tmp_V_68_fu_1530 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd68))) begin
        tmp_V_69_fu_1534 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd5))) begin
        tmp_V_6_fu_1282 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd69))) begin
        tmp_V_70_fu_1538 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd70))) begin
        tmp_V_71_fu_1542 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd71))) begin
        tmp_V_72_fu_1546 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd72))) begin
        tmp_V_73_fu_1550 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd73))) begin
        tmp_V_74_fu_1554 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd74))) begin
        tmp_V_75_fu_1558 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd75))) begin
        tmp_V_76_fu_1562 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd76))) begin
        tmp_V_77_fu_1566 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd77))) begin
        tmp_V_78_fu_1570 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd78))) begin
        tmp_V_79_fu_1574 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd6))) begin
        tmp_V_7_fu_1286 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd79))) begin
        tmp_V_80_fu_1578 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd80))) begin
        tmp_V_81_fu_1582 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd81))) begin
        tmp_V_82_fu_1586 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd82))) begin
        tmp_V_83_fu_1590 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd83))) begin
        tmp_V_84_fu_1594 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd84))) begin
        tmp_V_85_fu_1598 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd85))) begin
        tmp_V_86_fu_1602 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd86))) begin
        tmp_V_87_fu_1606 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd87))) begin
        tmp_V_88_fu_1610 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd88))) begin
        tmp_V_89_fu_1614 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd7))) begin
        tmp_V_8_fu_1290 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd89))) begin
        tmp_V_90_fu_1618 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd90))) begin
        tmp_V_91_fu_1622 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd91))) begin
        tmp_V_92_fu_1626 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd92))) begin
        tmp_V_93_fu_1630 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd93))) begin
        tmp_V_94_fu_1634 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd94))) begin
        tmp_V_95_fu_1638 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd95))) begin
        tmp_V_96_fu_1642 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd96))) begin
        tmp_V_97_fu_1646 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd97))) begin
        tmp_V_98_fu_1650 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd98))) begin
        tmp_V_99_fu_1654 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd8))) begin
        tmp_V_9_fu_1294 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_7683_p1 == 10'd0))) begin
        tmp_V_fu_1262 <= in_V_V_TDATA;
    end
end

always @ (*) begin
    if ((icmp_ln248_fu_4769_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_15104 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_sig_allocacmp_nf_0_load_1 = select_ln301_fu_10945_p3;
    end else begin
        ap_sig_allocacmp_nf_0_load_1 = nf_0_fu_3566;
    end
end

always @ (*) begin
    if (((icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op1183_read_state2 == 1'b1))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_15104 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_15104 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln248_fu_4769_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TDATA_blk_n = weight_V_V_TVALID;
    end else begin
        weight_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_4769_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TREADY = 1'b1;
    end else begin
        weight_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((icmp_ln248_fu_4769_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((icmp_ln248_fu_4769_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accu_0_0_V_fu_10765_p2 = ($signed(select_ln271_3_fu_10700_p3) + $signed(sext_ln700_1_fu_10761_p1));

assign accu_0_1_V_fu_10807_p2 = ($signed(select_ln271_2_fu_10693_p3) + $signed(sext_ln700_3_fu_10803_p1));

assign accu_0_2_V_fu_10849_p2 = ($signed(select_ln271_1_fu_10686_p3) + $signed(sext_ln700_5_fu_10845_p1));

assign accu_0_3_V_fu_10891_p2 = ($signed(select_ln271_fu_10679_p3) + $signed(sext_ln700_7_fu_10887_p1));

assign add_ln700_2_fu_10797_p2 = ($signed(sext_ln700_2_fu_10793_p1) + $signed(sext_ln170_1_fu_10780_p1));

assign add_ln700_4_fu_10839_p2 = ($signed(sext_ln700_4_fu_10835_p1) + $signed(sext_ln170_2_fu_10822_p1));

assign add_ln700_6_fu_10881_p2 = ($signed(sext_ln700_6_fu_10877_p1) + $signed(sext_ln170_3_fu_10864_p1));

assign add_ln700_fu_10755_p2 = ($signed(sext_ln700_fu_10751_p1) + $signed(sext_ln170_fu_10724_p1));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op1183_read_state2 == 1'b1)) | ((icmp_ln248_fu_4769_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op1183_read_state2 == 1'b1)) | ((icmp_ln248_fu_4769_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op1183_read_state2 == 1'b1)) | ((icmp_ln248_fu_4769_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op1183_read_state2 == 1'b1)) | ((icmp_ln248_fu_4769_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)));
end

always @ (*) begin
    ap_block_state3_io = ((icmp_ln289_reg_15104 == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_reg_pp0_iter0_act_m_val_V_reg_3600 = 'bx;

always @ (*) begin
    ap_predicate_op1183_read_state2 = ((icmp_ln252_fu_4784_p2 == 1'd1) & (icmp_ln248_fu_4769_p2 == 1'd0));
end

assign arg_V_read_assign_1_fu_10728_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_3600[7:4]}};

assign i_fu_4775_p2 = (i_0_reg_3589 + 21'd1);

assign icmp_ln248_fu_4769_p2 = ((i_0_reg_3589 == 21'd1843200) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_4784_p2 = ((ap_sig_allocacmp_nf_0_load_1 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln271_fu_10570_p2 = ((sf_1_fu_1258 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln289_fu_10656_p2 = ((sf_fu_10650_p2 == 32'd576) ? 1'b1 : 1'b0);

assign icmp_ln301_fu_10939_p2 = ((nf_fu_10933_p2 == 32'd32) ? 1'b1 : 1'b0);

assign inElem_V_1_fu_6525_p577 = sf_1_fu_1258[9:0];

assign mul_ln1352_1_fu_10745_p0 = sext_ln215_3_fu_10741_p1;

assign mul_ln1352_2_fu_10774_p0 = sext_ln215_1_fu_10714_p1;

assign mul_ln1352_3_fu_10787_p0 = sext_ln215_3_fu_10741_p1;

assign mul_ln1352_4_fu_10816_p0 = sext_ln215_1_fu_10714_p1;

assign mul_ln1352_5_fu_10829_p0 = sext_ln215_3_fu_10741_p1;

assign mul_ln1352_6_fu_10858_p0 = sext_ln215_1_fu_10714_p1;

assign mul_ln1352_7_fu_10871_p0 = sext_ln215_3_fu_10741_p1;

assign mul_ln1352_fu_10718_p0 = sext_ln215_1_fu_10714_p1;

assign nf_fu_10933_p2 = (nf_0_fu_3566 + 32'd1);

assign out_V_V_TDATA = {{{{accu_0_3_V_fu_10891_p2}, {accu_0_2_V_fu_10849_p2}}, {accu_0_1_V_fu_10807_p2}}, {accu_0_0_V_fu_10765_p2}};

assign select_ln271_1_fu_10686_p3 = ((icmp_ln271_reg_15056[0:0] === 1'b1) ? 24'd0 : accu_0_2_V_1_fu_1250);

assign select_ln271_2_fu_10693_p3 = ((icmp_ln271_reg_15056[0:0] === 1'b1) ? 24'd0 : accu_0_1_V_1_fu_1246);

assign select_ln271_3_fu_10700_p3 = ((icmp_ln271_reg_15056[0:0] === 1'b1) ? 24'd0 : accu_0_0_V_1_fu_1242);

assign select_ln271_fu_10679_p3 = ((icmp_ln271_reg_15056[0:0] === 1'b1) ? 24'd0 : accu_0_3_V_1_fu_1254);

assign select_ln301_fu_10945_p3 = ((icmp_ln301_fu_10939_p2[0:0] === 1'b1) ? 32'd0 : nf_fu_10933_p2);

assign sext_ln170_1_fu_10780_p1 = mul_ln1352_2_fu_10774_p2;

assign sext_ln170_2_fu_10822_p1 = mul_ln1352_4_fu_10816_p2;

assign sext_ln170_3_fu_10864_p1 = mul_ln1352_6_fu_10858_p2;

assign sext_ln170_fu_10724_p1 = mul_ln1352_fu_10718_p2;

assign sext_ln215_1_fu_10714_p1 = $signed(trunc_ln647_1_fu_10707_p1);

assign sext_ln215_3_fu_10741_p1 = $signed(arg_V_read_assign_1_fu_10728_p4);

assign sext_ln700_1_fu_10761_p1 = $signed(add_ln700_fu_10755_p2);

assign sext_ln700_2_fu_10793_p1 = mul_ln1352_3_fu_10787_p2;

assign sext_ln700_3_fu_10803_p1 = $signed(add_ln700_2_fu_10797_p2);

assign sext_ln700_4_fu_10835_p1 = mul_ln1352_5_fu_10829_p2;

assign sext_ln700_5_fu_10845_p1 = $signed(add_ln700_4_fu_10839_p2);

assign sext_ln700_6_fu_10877_p1 = mul_ln1352_7_fu_10871_p2;

assign sext_ln700_7_fu_10887_p1 = $signed(add_ln700_6_fu_10881_p2);

assign sext_ln700_fu_10751_p1 = mul_ln1352_1_fu_10745_p2;

assign sf_fu_10650_p2 = (32'd1 + sf_1_fu_1258);

assign trunc_ln321_fu_7683_p1 = sf_1_fu_1258[9:0];

assign trunc_ln647_1_fu_10707_p1 = ap_phi_reg_pp0_iter1_act_m_val_V_reg_3600[3:0];

assign trunc_ln647_fu_10576_p1 = weight_V_V_TDATA[3:0];

endmodule //StreamingFCLayer_Batch_0_Matrix_Vector_Activa
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActLf8.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActLf8_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActLf8_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActLf8(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActLf8_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActLf8_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActHfu.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActHfu_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActHfu_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActHfu(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActHfu_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActHfu_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcsc4.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcsc4_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 5;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcsc4_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcsc4(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd5;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcsc4_rom Thresholding_Batch_0_Thresholding_Batcsc4_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActOgC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActOgC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActOgC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActOgC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActOgC_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActOgC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc3C.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcc3C_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc3C_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcc3C(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcc3C_rom Thresholding_Batch_0_Thresholding_Batcc3C_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Acthbi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Acthbi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Acthbi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Acthbi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Acthbi_rom StreamingFCLayer_Batch_1_Matrix_Vector_Acthbi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_BatceOg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_BatceOg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_BatceOg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_BatceOg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_BatceOg_rom Thresholding_Batch_2_Thresholding_BatceOg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/6c99/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActPgM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActPgM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActPgM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActPgM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActPgM_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActPgM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8b1e/StreamingFIFO_5.v


module StreamingFIFO_5(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(16)
)
StreamingFIFO_5_StreamingFIFO_5
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/209a/hdl/mux.v

/*
 Copyright (c) 2020, Xilinx
 All rights reserved.

 Redistribution and use in source and binary forms, with or without
 modification, are permitted provided that the following conditions are met:

 * Redistributions of source code must retain the above copyright notice, this
   list of conditions and the following disclaimer.

 * Redistributions in binary form must reproduce the above copyright notice,
   this list of conditions and the following disclaimer in the documentation
   and/or other materials provided with the distribution.

 * Neither the name of FINN nor the names of its
   contributors may be used to endorse or promote products derived from
   this software without specific prior written permission.

 THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
 FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
 SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
 CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
 OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

module mux
#(
    parameter NINPUTS = 1,
	parameter WIDTH = 16
)
(
	input [NINPUTS*WIDTH-1:0] in,
	output [WIDTH-1:0] out,
	input [$clog2(NINPUTS)-1:0] sel
);

assign out = in >> (sel*WIDTH);

endmodule//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbil.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbil_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbil_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbil(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbil_rom Thresholding_Batch_0_Thresholding_Batcbil_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActqcK.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActqcK_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActqcK_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActqcK(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActqcK_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActqcK_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActZio.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActZio_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActZio_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActZio(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActZio_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActZio_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbHp.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcbHp_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbHp_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcbHp(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcbHp_rom Thresholding_Batch_0_Thresholding_BatcbHp_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcckv.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcckv_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcckv_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcckv(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcckv_rom Thresholding_Batch_0_Thresholding_Batcckv_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_Batch_2.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="Thresholding_Batch_2_Thresholding_Batch_2,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.733750,HLS_SYN_LAT=50182,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=578,HLS_SYN_LUT=895,HLS_VERSION=2020_1_1}" *)

module Thresholding_Batch_2_Thresholding_Batch_2 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_Thresholding_Batch_fu_60_ap_start;
wire    grp_Thresholding_Batch_fu_60_ap_done;
wire    grp_Thresholding_Batch_fu_60_ap_idle;
wire    grp_Thresholding_Batch_fu_60_ap_ready;
wire    grp_Thresholding_Batch_fu_60_in_V_V_TREADY;
wire   [7:0] grp_Thresholding_Batch_fu_60_out_V_V_TDATA;
wire    grp_Thresholding_Batch_fu_60_out_V_V_TVALID;
wire    grp_Thresholding_Batch_fu_60_out_V_V_TREADY;
reg    grp_Thresholding_Batch_fu_60_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [15:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_Thresholding_Batch_fu_60_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

Thresholding_Batch_2_Thresholding_Batch grp_Thresholding_Batch_fu_60(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_Thresholding_Batch_fu_60_ap_start),
    .ap_done(grp_Thresholding_Batch_fu_60_ap_done),
    .ap_idle(grp_Thresholding_Batch_fu_60_ap_idle),
    .ap_ready(grp_Thresholding_Batch_fu_60_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_Thresholding_Batch_fu_60_in_V_V_TREADY),
    .out_V_V_TDATA(grp_Thresholding_Batch_fu_60_out_V_V_TDATA),
    .out_V_V_TVALID(grp_Thresholding_Batch_fu_60_out_V_V_TVALID),
    .out_V_V_TREADY(grp_Thresholding_Batch_fu_60_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_Thresholding_Batch_fu_60_out_V_V_TDATA),
    .vld_in(grp_Thresholding_Batch_fu_60_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_Thresholding_Batch_fu_60_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_Thresholding_Batch_fu_60_ap_start_reg <= 1'b1;
        end else if ((grp_Thresholding_Batch_fu_60_ap_ready == 1'b1)) begin
            grp_Thresholding_Batch_fu_60_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_Thresholding_Batch_fu_60_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_Thresholding_Batch_fu_60_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((1'b1 == ap_CS_fsm_state4) & (regslice_both_out_V_V_U_apdone_blk == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_Thresholding_Batch_fu_60_ap_start = grp_Thresholding_Batch_fu_60_ap_start_reg;

assign grp_Thresholding_Batch_fu_60_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //Thresholding_Batch_2_Thresholding_Batch_2
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActLf8.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActLf8_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActLf8_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActLf8(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActLf8_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActLf8_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Act1iI.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Act1iI_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Act1iI_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Act1iI(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Act1iI_rom StreamingFCLayer_Batch_1_Matrix_Vector_Act1iI_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdaE.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcdaE_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdaE_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcdaE(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcdaE_rom Thresholding_Batch_0_Thresholding_BatcdaE_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActxdS.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActxdS_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActxdS_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActxdS(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActxdS_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActxdS_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8799/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccpw.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccpw_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccpw_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccpw(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccpw_rom Thresholding_Batch_0_Thresholding_Batccpw_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_StreamingFCLayer_5jm.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module StreamingFCLayer_Batch_2_StreamingFCLayer_5jm #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH       = 32,
    din5_WIDTH       = 32,
    din6_WIDTH       = 32,
    din7_WIDTH       = 32,
    din8_WIDTH       = 32,
    din9_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [23 : 0]     din0,
    input  [23 : 0]     din1,
    input  [23 : 0]     din2,
    input  [23 : 0]     din3,
    input  [23 : 0]     din4,
    input  [23 : 0]     din5,
    input  [23 : 0]     din6,
    input  [23 : 0]     din7,
    input  [23 : 0]     din8,
    input  [3 : 0]    din9,
    output [23 : 0]   dout);

// puts internal signals
wire [3 : 0]     sel;
// level 1 signals
wire [23 : 0]         mux_1_0;
wire [23 : 0]         mux_1_1;
wire [23 : 0]         mux_1_2;
wire [23 : 0]         mux_1_3;
wire [23 : 0]         mux_1_4;
// level 2 signals
wire [23 : 0]         mux_2_0;
wire [23 : 0]         mux_2_1;
wire [23 : 0]         mux_2_2;
// level 3 signals
wire [23 : 0]         mux_3_0;
wire [23 : 0]         mux_3_1;
// level 4 signals
wire [23 : 0]         mux_4_0;

assign sel = din9;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;
assign mux_1_2 = (sel[0] == 0)? din4 : din5;
assign mux_1_3 = (sel[0] == 0)? din6 : din7;
assign mux_1_4 = din8;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;
assign mux_2_1 = (sel[1] == 0)? mux_1_2 : mux_1_3;
assign mux_2_2 = mux_1_4;

// Generate level 3 logic
assign mux_3_0 = (sel[2] == 0)? mux_2_0 : mux_2_1;
assign mux_3_1 = mux_2_2;

// Generate level 4 logic
assign mux_4_0 = (sel[3] == 0)? mux_3_0 : mux_3_1;

// output logic
assign dout = mux_4_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actbkb_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actbkb_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actbkb(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actbkb_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actbkb_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatckbM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatckbM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 4;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatckbM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatckbM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd4;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatckbM_rom Thresholding_Batch_0_Thresholding_BatckbM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbdk.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbdk_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbdk_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbdk(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbdk_rom Thresholding_Batch_0_Thresholding_Batcbdk_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_4_wstrm_0/synth/finn_design_StreamingFCLayer_Batch_4_wstrm_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:user:memstream:1.0
// IP Revision: 5

(* X_CORE_INFO = "memstream,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_4_wstrm_0,memstream,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_4_wstrm_0,memstream,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=user,x_ipName=memstream,x_ipVersion=1.0,x_ipCoreRevision=5,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED,CONFIG_EN=true,NSTREAMS=1,MEM_DEPTH=8192,MEM_WIDTH=128,MEM_INIT=/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/,RAM_STYLE=auto,STRM0_WIDTH=128,STRM1_WIDTH=32,STRM2_WIDTH=32,STRM3_WIDTH=32,STRM4_WIDTH=32,STRM5_WIDTH=32,ST\
RM0_DEPTH=8192,STRM1_DEPTH=2304,STRM2_DEPTH=2304,STRM3_DEPTH=2304,STRM4_DEPTH=2304,STRM5_DEPTH=2304,STRM0_OFFSET=0,STRM1_OFFSET=2304,STRM2_OFFSET=4608,STRM3_OFFSET=6912,STRM4_OFFSET=9216,STRM5_OFFSET=11520,AXILITE_ADDR_WIDTH=17}" *)
(* IP_DEFINITION_SOURCE = "package_project" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_4_wstrm_0 (
  aclk,
  aresetn,
  awready,
  awvalid,
  awaddr,
  awprot,
  wready,
  wvalid,
  wdata,
  wstrb,
  bready,
  bvalid,
  bresp,
  arready,
  arvalid,
  araddr,
  arprot,
  rready,
  rvalid,
  rresp,
  rdata,
  m_axis_0_tready,
  m_axis_0_tvalid,
  m_axis_0_tdata
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aclk, ASSOCIATED_BUSIF m_axis_0:m_axis_1:m_axis_2:m_axis_3:m_axis_4:m_axis_5:s_axilite, ASSOCIATED_RESET aresetn, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 aclk CLK" *)
input wire aclk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aresetn, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 aresetn RST" *)
input wire aresetn;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWREADY" *)
output wire awready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWVALID" *)
input wire awvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWADDR" *)
input wire [16 : 0] awaddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWPROT" *)
input wire [2 : 0] awprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WREADY" *)
output wire wready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WVALID" *)
input wire wvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WDATA" *)
input wire [31 : 0] wdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WSTRB" *)
input wire [3 : 0] wstrb;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BREADY" *)
input wire bready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BVALID" *)
output wire bvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BRESP" *)
output wire [1 : 0] bresp;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARREADY" *)
output wire arready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARVALID" *)
input wire arvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARADDR" *)
input wire [16 : 0] araddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARPROT" *)
input wire [2 : 0] arprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RREADY" *)
input wire rready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RVALID" *)
output wire rvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RRESP" *)
output wire [1 : 0] rresp;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axilite, DATA_WIDTH 32, PROTOCOL AXI4LITE, FREQ_HZ 100000000.000000, ID_WIDTH 0, ADDR_WIDTH 17, AWUSER_WIDTH 0, ARUSER_WIDTH 0, WUSER_WIDTH 0, RUSER_WIDTH 0, BUSER_WIDTH 0, READ_WRITE_MODE READ_WRITE, HAS_BURST 0, HAS_LOCK 0, HAS_PROT 1, HAS_CACHE 0, HAS_QOS 0, HAS_REGION 0, HAS_WSTRB 1, HAS_BRESP 1, HAS_RRESP 1, SUPPORTS_NARROW_BURST 0, NUM_READ_OUTSTANDING 1, NUM_WRITE_OUTSTANDING 1, MAX_BURST_LENGTH 1, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, NUM_READ_THREADS 1, NUM_W\
RITE_THREADS 1, RUSER_BITS_PER_BYTE 0, WUSER_BITS_PER_BYTE 0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RDATA" *)
output wire [31 : 0] rdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TREADY" *)
input wire m_axis_0_tready;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TVALID" *)
output wire m_axis_0_tvalid;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME m_axis_0, TDATA_NUM_BYTES 16, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TDATA" *)
output wire [127 : 0] m_axis_0_tdata;

  memstream #(
    .CONFIG_EN(1'B1),
    .NSTREAMS(1),
    .MEM_DEPTH(8192),
    .MEM_WIDTH(128),
    .MEM_INIT("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/"),
    .RAM_STYLE("auto"),
    .STRM0_WIDTH(128),
    .STRM1_WIDTH(32),
    .STRM2_WIDTH(32),
    .STRM3_WIDTH(32),
    .STRM4_WIDTH(32),
    .STRM5_WIDTH(32),
    .STRM0_DEPTH(8192),
    .STRM1_DEPTH(2304),
    .STRM2_DEPTH(2304),
    .STRM3_DEPTH(2304),
    .STRM4_DEPTH(2304),
    .STRM5_DEPTH(2304),
    .STRM0_OFFSET(0),
    .STRM1_OFFSET(2304),
    .STRM2_OFFSET(4608),
    .STRM3_OFFSET(6912),
    .STRM4_OFFSET(9216),
    .STRM5_OFFSET(11520),
    .AXILITE_ADDR_WIDTH(17)
  ) inst (
    .aclk(aclk),
    .aresetn(aresetn),
    .awready(awready),
    .awvalid(awvalid),
    .awaddr(awaddr),
    .awprot(awprot),
    .wready(wready),
    .wvalid(wvalid),
    .wdata(wdata),
    .wstrb(wstrb),
    .bready(bready),
    .bvalid(bvalid),
    .bresp(bresp),
    .arready(arready),
    .arvalid(arvalid),
    .araddr(araddr),
    .arprot(arprot),
    .rready(rready),
    .rvalid(rvalid),
    .rresp(rresp),
    .rdata(rdata),
    .m_axis_0_afull(1'B0),
    .m_axis_0_tready(m_axis_0_tready),
    .m_axis_0_tvalid(m_axis_0_tvalid),
    .m_axis_0_tdata(m_axis_0_tdata),
    .m_axis_1_afull(1'B0),
    .m_axis_1_tready(1'B1),
    .m_axis_1_tvalid(),
    .m_axis_1_tdata(),
    .m_axis_2_afull(1'B0),
    .m_axis_2_tready(1'B1),
    .m_axis_2_tvalid(),
    .m_axis_2_tdata(),
    .m_axis_3_afull(1'B0),
    .m_axis_3_tready(1'B1),
    .m_axis_3_tvalid(),
    .m_axis_3_tdata(),
    .m_axis_4_afull(1'B0),
    .m_axis_4_tready(1'B1),
    .m_axis_4_tvalid(),
    .m_axis_4_tdata(),
    .m_axis_5_afull(1'B0),
    .m_axis_5_tready(1'B1),
    .m_axis_5_tvalid(),
    .m_axis_5_tdata()
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actudo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actudo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actudo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actudo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actudo_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actudo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActkbM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActkbM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActkbM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActkbM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActkbM_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActkbM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActFfa.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActFfa_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActFfa_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActFfa(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActFfa_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActFfa_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActThq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActThq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActThq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActThq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActThq_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActThq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActVhK.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActVhK_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActVhK_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActVhK(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActVhK_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActVhK_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Act4jc.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Act4jc_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Act4jc_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Act4jc(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Act4jc_rom StreamingFCLayer_Batch_4_Matrix_Vector_Act4jc_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcczy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcczy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcczy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcczy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcczy_rom Thresholding_Batch_0_Thresholding_Batcczy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Act4jc.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Act4jc_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Act4jc_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Act4jc(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Act4jc_rom StreamingFCLayer_Batch_1_Matrix_Vector_Act4jc_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccZC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccZC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccZC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccZC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccZC_rom Thresholding_Batch_0_Thresholding_BatccZC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_3_0/synth/finn_design_StreamingFIFO_3_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_3:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_3,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_3_0,StreamingFIFO_3,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_3_0,StreamingFIFO_3,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_3,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_3_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [7 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_3 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_Batch_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="Thresholding_Batch_1_Thresholding_Batch_1,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.079000,HLS_SYN_LAT=12806,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=629,HLS_SYN_LUT=1179,HLS_VERSION=2020_1_1}" *)

module Thresholding_Batch_1_Thresholding_Batch_1 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [23:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_Thresholding_Batch_fu_60_ap_start;
wire    grp_Thresholding_Batch_fu_60_ap_done;
wire    grp_Thresholding_Batch_fu_60_ap_idle;
wire    grp_Thresholding_Batch_fu_60_ap_ready;
wire    grp_Thresholding_Batch_fu_60_in_V_V_TREADY;
wire   [7:0] grp_Thresholding_Batch_fu_60_out_V_V_TDATA;
wire    grp_Thresholding_Batch_fu_60_out_V_V_TVALID;
wire    grp_Thresholding_Batch_fu_60_out_V_V_TREADY;
reg    grp_Thresholding_Batch_fu_60_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [23:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_Thresholding_Batch_fu_60_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

Thresholding_Batch_1_Thresholding_Batch grp_Thresholding_Batch_fu_60(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_Thresholding_Batch_fu_60_ap_start),
    .ap_done(grp_Thresholding_Batch_fu_60_ap_done),
    .ap_idle(grp_Thresholding_Batch_fu_60_ap_idle),
    .ap_ready(grp_Thresholding_Batch_fu_60_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_Thresholding_Batch_fu_60_in_V_V_TREADY),
    .out_V_V_TDATA(grp_Thresholding_Batch_fu_60_out_V_V_TDATA),
    .out_V_V_TVALID(grp_Thresholding_Batch_fu_60_out_V_V_TVALID),
    .out_V_V_TREADY(grp_Thresholding_Batch_fu_60_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 24 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_Thresholding_Batch_fu_60_out_V_V_TDATA),
    .vld_in(grp_Thresholding_Batch_fu_60_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_Thresholding_Batch_fu_60_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_Thresholding_Batch_fu_60_ap_start_reg <= 1'b1;
        end else if ((grp_Thresholding_Batch_fu_60_ap_ready == 1'b1)) begin
            grp_Thresholding_Batch_fu_60_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_Thresholding_Batch_fu_60_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_Thresholding_Batch_fu_60_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((1'b1 == ap_CS_fsm_state4) & (regslice_both_out_V_V_U_apdone_blk == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_Thresholding_Batch_fu_60_ap_start = grp_Thresholding_Batch_fu_60_ap_start_reg;

assign grp_Thresholding_Batch_fu_60_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //Thresholding_Batch_1_Thresholding_Batch_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcUhA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcUhA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcUhA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcUhA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcUhA_rom Thresholding_Batch_0_Thresholding_BatcUhA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingDataWidthConverter_Batch_2_0/synth/finn_design_StreamingDataWidthConverter_Batch_2_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingDataWidthConverter_Batch_2:1.0
// IP Revision: 2101301322

(* X_CORE_INFO = "StreamingDataWidthConverter_Batch_2_StreamingDataWidthConverter_Batch_2,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingDataWidthConverter_Batch_2_0,StreamingDataWidthConverter_Batch_2_StreamingDataWidthConverter_Batch_2,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingDataWidthConverter_Batch_2_0,StreamingDataWidthConverter_Batch_2_StreamingDataWidthConverter_Batch_2,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingDataWidthConverter_Batch_2,x_ipVersion=1.0,x_ipCoreRevision=2101301322,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingDataWidthConverter_Batch_2_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 4, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [31 : 0] out_V_V_TDATA;

  StreamingDataWidthConverter_Batch_2_StreamingDataWidthConverter_Batch_2 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actsc4.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actsc4_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actsc4_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actsc4(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actsc4_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actsc4_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Act2iS.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Act2iS_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Act2iS_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Act2iS(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Act2iS_rom StreamingFCLayer_Batch_2_Matrix_Vector_Act2iS_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actzec.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actzec_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actzec_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actzec(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actzec_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actzec_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/be37/StreamingFIFO_13.v


module StreamingFIFO_13(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [31:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(32)
)
StreamingFIFO_13_StreamingFIFO_13
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actncg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actncg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actncg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actncg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actncg_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actncg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/e03c/hdl/verilog/ConvolutionInputGenerator_3_ConvolutionInputGene_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module ConvolutionInputGenerator_3_ConvolutionInputGene_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [31:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln197_fu_374_p2;
wire   [0:0] icmp_ln199_fu_396_p2;
wire   [0:0] and_ln245_fu_606_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln199_reg_893;
reg   [0:0] icmp_ln215_reg_897;
reg   [15:0] i_0_0_reg_277;
reg    ap_predicate_op119_read_state2;
reg    ap_predicate_op162_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_predicate_op205_write_state3;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [15:0] add_ln197_fu_380_p2;
wire   [0:0] icmp_ln215_fu_405_p2;
wire   [1:0] add_ln221_fu_479_p2;
reg   [1:0] add_ln221_reg_901;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
wire   [7:0] inputBuf_0_V_address0;
reg    inputBuf_0_V_ce0;
wire   [31:0] inputBuf_0_V_q0;
reg   [7:0] inputBuf_0_V_address1;
reg    inputBuf_0_V_ce1;
reg    inputBuf_0_V_we1;
wire   [7:0] inputBuf_1_V_address0;
reg    inputBuf_1_V_ce0;
wire   [31:0] inputBuf_1_V_q0;
reg   [7:0] inputBuf_1_V_address1;
reg    inputBuf_1_V_ce1;
reg    inputBuf_1_V_we1;
wire   [7:0] inputBuf_2_V_address0;
reg    inputBuf_2_V_ce0;
wire   [31:0] inputBuf_2_V_q0;
reg   [7:0] inputBuf_2_V_address1;
reg    inputBuf_2_V_ce1;
reg    inputBuf_2_V_we1;
wire   [7:0] inputBuf_3_V_address0;
reg    inputBuf_3_V_ce0;
wire   [31:0] inputBuf_3_V_q0;
reg   [7:0] inputBuf_3_V_address1;
reg    inputBuf_3_V_ce1;
reg    inputBuf_3_V_we1;
wire   [63:0] zext_ln221_fu_465_p1;
wire   [63:0] zext_ln248_fu_612_p1;
wire   [63:0] zext_ln202_fu_724_p1;
reg   [31:0] ofm_y_1_0_fu_84;
wire   [31:0] select_ln236_1_fu_573_p3;
wire   [0:0] icmp_ln224_fu_491_p2;
wire   [0:0] icmp_ln227_fu_508_p2;
wire   [0:0] icmp_ln230_fu_519_p2;
wire   [0:0] icmp_ln233_fu_539_p2;
reg   [31:0] ofm_x_1_0_fu_88;
wire   [31:0] add_ln232_fu_533_p2;
reg   [31:0] k_y_1_0_fu_92;
wire   [31:0] add_ln216_fu_427_p2;
reg   [31:0] inp_15_0_fu_96;
wire   [31:0] select_ln236_fu_565_p3;
wire   [31:0] add_ln204_fu_736_p2;
reg   [31:0] k_x_1_0_fu_100;
wire   [31:0] add_ln226_fu_502_p2;
reg   [31:0] count_simd_1_0_fu_104;
wire   [31:0] add_ln223_fu_485_p2;
reg   [31:0] read_block_1_0_fu_108;
wire   [31:0] zext_ln252_fu_677_p1;
wire   [31:0] add_ln211_fu_772_p2;
wire   [0:0] icmp_ln205_fu_348_p2;
reg   [31:0] current_block_write_s_fu_112;
wire   [31:0] select_ln252_fu_653_p3;
wire   [31:0] select_ln208_fu_764_p3;
reg   [31:0] current_line_1_0_fu_116;
wire   [31:0] select_ln252_1_fu_661_p3;
wire   [31:0] grp_fu_336_p2;
reg   [31:0] counter_internal_blo_fu_120;
wire   [31:0] select_ln264_fu_711_p3;
wire   [31:0] tmp_V_1_fu_788_p6;
reg    ap_block_pp0_stage0_01001;
wire   [1:0] trunc_ln321_1_fu_620_p1;
wire   [1:0] trunc_ln321_fu_732_p1;
wire   [28:0] trunc_ln220_1_fu_441_p1;
wire   [28:0] trunc_ln220_fu_437_p1;
wire   [28:0] add_ln220_fu_445_p2;
wire   [31:0] shl_ln_fu_451_p3;
wire   [31:0] add_ln220_1_fu_459_p2;
wire   [1:0] trunc_ln216_1_fu_433_p1;
wire   [1:0] add_ln221_1_fu_473_p2;
wire   [1:0] trunc_ln216_fu_423_p1;
wire   [31:0] add_ln235_fu_553_p2;
wire   [0:0] icmp_ln236_fu_559_p2;
wire   [0:0] icmp_ln245_fu_594_p2;
wire   [0:0] icmp_ln245_1_fu_600_p2;
wire   [4:0] trunc_ln197_fu_392_p1;
wire   [31:0] add_ln256_fu_633_p2;
wire   [0:0] icmp_ln257_fu_639_p2;
wire   [0:0] icmp_ln252_fu_342_p2;
wire   [31:0] select_ln257_fu_645_p3;
wire   [4:0] add_ln256_1_fu_627_p2;
wire   [4:0] select_ln252_2_fu_669_p3;
wire   [31:0] add_ln263_fu_699_p2;
wire   [0:0] icmp_ln264_fu_705_p2;
wire   [31:0] add_ln207_fu_752_p2;
wire   [0:0] icmp_ln208_fu_758_p2;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_block_pp0;
reg    ap_predicate_op127_store_state2;
reg    ap_enable_operation_127;
reg    ap_enable_state2_pp0_iter0_stage0;
reg    ap_predicate_op69_load_state2;
reg    ap_enable_operation_69;
reg    ap_predicate_op202_load_state3;
reg    ap_enable_operation_202;
reg    ap_enable_state3_pp0_iter1_stage0;
reg    ap_predicate_op170_store_state2;
reg    ap_enable_operation_170;
reg    ap_predicate_op129_store_state2;
reg    ap_enable_operation_129;
reg    ap_predicate_op67_load_state2;
reg    ap_enable_operation_67;
reg    ap_predicate_op201_load_state3;
reg    ap_enable_operation_201;
reg    ap_predicate_op172_store_state2;
reg    ap_enable_operation_172;
reg    ap_predicate_op131_store_state2;
reg    ap_enable_operation_131;
reg    ap_predicate_op65_load_state2;
reg    ap_enable_operation_65;
reg    ap_predicate_op200_load_state3;
reg    ap_enable_operation_200;
reg    ap_predicate_op174_store_state2;
reg    ap_enable_operation_174;
reg    ap_predicate_op133_store_state2;
reg    ap_enable_operation_133;
reg    ap_predicate_op71_load_state2;
reg    ap_enable_operation_71;
reg    ap_predicate_op203_load_state3;
reg    ap_enable_operation_203;
reg    ap_predicate_op176_store_state2;
reg    ap_enable_operation_176;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_660;
reg    ap_condition_230;
reg    ap_condition_666;
reg    ap_condition_670;
reg    ap_condition_674;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

ConvolutionInputGenerator_3_ConvolutionInputGbkb #(
    .DataWidth( 32 ),
    .AddressRange( 240 ),
    .AddressWidth( 8 ))
inputBuf_0_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_0_V_address0),
    .ce0(inputBuf_0_V_ce0),
    .q0(inputBuf_0_V_q0),
    .address1(inputBuf_0_V_address1),
    .ce1(inputBuf_0_V_ce1),
    .we1(inputBuf_0_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_3_ConvolutionInputGbkb #(
    .DataWidth( 32 ),
    .AddressRange( 240 ),
    .AddressWidth( 8 ))
inputBuf_1_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_1_V_address0),
    .ce0(inputBuf_1_V_ce0),
    .q0(inputBuf_1_V_q0),
    .address1(inputBuf_1_V_address1),
    .ce1(inputBuf_1_V_ce1),
    .we1(inputBuf_1_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_3_ConvolutionInputGbkb #(
    .DataWidth( 32 ),
    .AddressRange( 240 ),
    .AddressWidth( 8 ))
inputBuf_2_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_2_V_address0),
    .ce0(inputBuf_2_V_ce0),
    .q0(inputBuf_2_V_q0),
    .address1(inputBuf_2_V_address1),
    .ce1(inputBuf_2_V_ce1),
    .we1(inputBuf_2_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_3_ConvolutionInputGbkb #(
    .DataWidth( 32 ),
    .AddressRange( 240 ),
    .AddressWidth( 8 ))
inputBuf_3_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_3_V_address0),
    .ce0(inputBuf_3_V_ce0),
    .q0(inputBuf_3_V_q0),
    .address1(inputBuf_3_V_address1),
    .ce1(inputBuf_3_V_ce1),
    .we1(inputBuf_3_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_3_ConvolutionInputGfYi #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
ConvolutionInputGfYi_U1(
    .din0(inputBuf_0_V_q0),
    .din1(inputBuf_1_V_q0),
    .din2(inputBuf_2_V_q0),
    .din3(inputBuf_3_V_q0),
    .din4(add_ln221_reg_901),
    .dout(tmp_V_1_fu_788_p6)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln224_fu_491_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        count_simd_1_0_fu_104 <= add_ln223_fu_485_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln227_fu_508_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln230_fu_519_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln233_fu_539_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln233_fu_539_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        count_simd_1_0_fu_104 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        counter_internal_blo_fu_120 <= select_ln264_fu_711_p3;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_348_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        counter_internal_blo_fu_120 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_348_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_block_write_s_fu_112 <= select_ln208_fu_764_p3;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_block_write_s_fu_112 <= select_ln252_fu_653_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        current_block_write_s_fu_112 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln205_fu_348_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_line_1_0_fu_116 <= grp_fu_336_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_line_1_0_fu_116 <= select_ln252_1_fu_661_p3;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_348_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        current_line_1_0_fu_116 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_0_reg_277 <= 16'd0;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_0_reg_277 <= add_ln197_fu_380_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inp_15_0_fu_96 <= add_ln204_fu_736_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln233_fu_539_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inp_15_0_fu_96 <= select_ln236_fu_565_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        inp_15_0_fu_96 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln227_fu_508_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        k_x_1_0_fu_100 <= add_ln226_fu_502_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln230_fu_519_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln233_fu_539_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln233_fu_539_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        k_x_1_0_fu_100 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln230_fu_519_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        k_y_1_0_fu_92 <= add_ln216_fu_427_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        k_y_1_0_fu_92 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln233_fu_539_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ofm_x_1_0_fu_88 <= add_ln232_fu_533_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln233_fu_539_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ofm_x_1_0_fu_88 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln233_fu_539_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ofm_y_1_0_fu_84 <= select_ln236_1_fu_573_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        ofm_y_1_0_fu_84 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_348_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        read_block_1_0_fu_108 <= add_ln211_fu_772_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        read_block_1_0_fu_108 <= zext_ln252_fu_677_p1;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        read_block_1_0_fu_108 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln221_reg_901 <= add_ln221_fu_479_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln197_fu_374_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln199_reg_893 <= icmp_ln199_fu_396_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln215_reg_897 <= icmp_ln215_fu_405_p2;
    end
end

always @ (*) begin
    if ((icmp_ln197_fu_374_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op119_read_state2 == 1'b1)))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_396_p2 == 1'd1) & (trunc_ln321_fu_732_p1 == 2'd0))) begin
            inputBuf_0_V_address1 = zext_ln202_fu_724_p1;
        end else if ((1'b1 == ap_condition_660)) begin
            inputBuf_0_V_address1 = zext_ln248_fu_612_p1;
        end else begin
            inputBuf_0_V_address1 = 'bx;
        end
    end else begin
        inputBuf_0_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_0_V_ce0 = 1'b1;
    end else begin
        inputBuf_0_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_0_V_ce1 = 1'b1;
    end else begin
        inputBuf_0_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_0_V_we1 = 1'b1;
    end else begin
        inputBuf_0_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_396_p2 == 1'd1) & (trunc_ln321_fu_732_p1 == 2'd1))) begin
            inputBuf_1_V_address1 = zext_ln202_fu_724_p1;
        end else if ((1'b1 == ap_condition_666)) begin
            inputBuf_1_V_address1 = zext_ln248_fu_612_p1;
        end else begin
            inputBuf_1_V_address1 = 'bx;
        end
    end else begin
        inputBuf_1_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_1_V_ce0 = 1'b1;
    end else begin
        inputBuf_1_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_1_V_ce1 = 1'b1;
    end else begin
        inputBuf_1_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_1_V_we1 = 1'b1;
    end else begin
        inputBuf_1_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_396_p2 == 1'd1) & (trunc_ln321_fu_732_p1 == 2'd2))) begin
            inputBuf_2_V_address1 = zext_ln202_fu_724_p1;
        end else if ((1'b1 == ap_condition_670)) begin
            inputBuf_2_V_address1 = zext_ln248_fu_612_p1;
        end else begin
            inputBuf_2_V_address1 = 'bx;
        end
    end else begin
        inputBuf_2_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_2_V_ce0 = 1'b1;
    end else begin
        inputBuf_2_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_2_V_ce1 = 1'b1;
    end else begin
        inputBuf_2_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_2_V_we1 = 1'b1;
    end else begin
        inputBuf_2_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_396_p2 == 1'd1) & (trunc_ln321_fu_732_p1 == 2'd3))) begin
            inputBuf_3_V_address1 = zext_ln202_fu_724_p1;
        end else if ((1'b1 == ap_condition_674)) begin
            inputBuf_3_V_address1 = zext_ln248_fu_612_p1;
        end else begin
            inputBuf_3_V_address1 = 'bx;
        end
    end else begin
        inputBuf_3_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_3_V_ce0 = 1'b1;
    end else begin
        inputBuf_3_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_3_V_ce1 = 1'b1;
    end else begin
        inputBuf_3_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_3_V_we1 = 1'b1;
    end else begin
        inputBuf_3_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op205_write_state3 == 1'b1))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((icmp_ln197_fu_374_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((icmp_ln197_fu_374_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln197_fu_380_p2 = (i_0_0_reg_277 + 16'd1);

assign add_ln204_fu_736_p2 = (inp_15_0_fu_96 + 32'd1);

assign add_ln207_fu_752_p2 = (current_block_write_s_fu_112 + 32'd1);

assign add_ln211_fu_772_p2 = (read_block_1_0_fu_108 + 32'd1);

assign add_ln216_fu_427_p2 = (32'd1 + k_y_1_0_fu_92);

assign add_ln220_1_fu_459_p2 = (shl_ln_fu_451_p3 + count_simd_1_0_fu_104);

assign add_ln220_fu_445_p2 = (trunc_ln220_1_fu_441_p1 + trunc_ln220_fu_437_p1);

assign add_ln221_1_fu_473_p2 = (2'd1 + trunc_ln216_1_fu_433_p1);

assign add_ln221_fu_479_p2 = (add_ln221_1_fu_473_p2 + trunc_ln216_fu_423_p1);

assign add_ln223_fu_485_p2 = (32'd1 + count_simd_1_0_fu_104);

assign add_ln226_fu_502_p2 = (k_x_1_0_fu_100 + 32'd1);

assign add_ln232_fu_533_p2 = (ofm_x_1_0_fu_88 + 32'd1);

assign add_ln235_fu_553_p2 = (ofm_y_1_0_fu_84 + 32'd1);

assign add_ln256_1_fu_627_p2 = (trunc_ln197_fu_392_p1 + 5'd1);

assign add_ln256_fu_633_p2 = (current_block_write_s_fu_112 + 32'd1);

assign add_ln263_fu_699_p2 = (counter_internal_blo_fu_120 + 32'd1);

assign and_ln245_fu_606_p2 = (icmp_ln245_fu_594_p2 & icmp_ln245_1_fu_600_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

always @ (*) begin
    ap_block_pp0 = ((ap_ST_fsm_pp0_stage0 == ap_CS_fsm) & (1'b1 == ap_block_pp0_stage0_subdone));
end

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1)));
end

always @ (*) begin
    ap_block_state3_io = ((out_V_V_TREADY == 1'b0) & (ap_predicate_op205_write_state3 == 1'b1));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_230 = ((icmp_ln197_fu_374_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_condition_660 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd0));
end

always @ (*) begin
    ap_condition_666 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd1));
end

always @ (*) begin
    ap_condition_670 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd2));
end

always @ (*) begin
    ap_condition_674 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd3));
end

always @ (*) begin
    ap_enable_operation_127 = (ap_predicate_op127_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_129 = (ap_predicate_op129_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_131 = (ap_predicate_op131_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_133 = (ap_predicate_op133_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_170 = (ap_predicate_op170_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_172 = (ap_predicate_op172_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_174 = (ap_predicate_op174_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_176 = (ap_predicate_op176_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_200 = (ap_predicate_op200_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_201 = (ap_predicate_op201_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_202 = (ap_predicate_op202_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_203 = (ap_predicate_op203_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_65 = (ap_predicate_op65_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_67 = (ap_predicate_op67_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_69 = (ap_predicate_op69_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_71 = (ap_predicate_op71_load_state2 == 1'b1);
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

always @ (*) begin
    ap_enable_state2_pp0_iter0_stage0 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_enable_state3_pp0_iter1_stage0 = ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_predicate_op119_read_state2 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op127_store_state2 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd2));
end

always @ (*) begin
    ap_predicate_op129_store_state2 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd1));
end

always @ (*) begin
    ap_predicate_op131_store_state2 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd0));
end

always @ (*) begin
    ap_predicate_op133_store_state2 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd3));
end

always @ (*) begin
    ap_predicate_op162_read_state2 = ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op170_store_state2 = ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd2));
end

always @ (*) begin
    ap_predicate_op172_store_state2 = ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd1));
end

always @ (*) begin
    ap_predicate_op174_store_state2 = ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd0));
end

always @ (*) begin
    ap_predicate_op176_store_state2 = ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd3));
end

always @ (*) begin
    ap_predicate_op200_load_state3 = ((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0));
end

always @ (*) begin
    ap_predicate_op201_load_state3 = ((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0));
end

always @ (*) begin
    ap_predicate_op202_load_state3 = ((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0));
end

always @ (*) begin
    ap_predicate_op203_load_state3 = ((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0));
end

always @ (*) begin
    ap_predicate_op205_write_state3 = ((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0));
end

always @ (*) begin
    ap_predicate_op65_load_state2 = ((icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op67_load_state2 = ((icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op69_load_state2 = ((icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op71_load_state2 = ((icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0));
end

assign grp_fu_336_p2 = (current_line_1_0_fu_116 + 32'd1);

assign icmp_ln197_fu_374_p2 = ((i_0_0_reg_277 == 16'd57168) ? 1'b1 : 1'b0);

assign icmp_ln199_fu_396_p2 = ((inp_15_0_fu_96 < 32'd720) ? 1'b1 : 1'b0);

assign icmp_ln205_fu_348_p2 = ((grp_fu_336_p2 == 32'd240) ? 1'b1 : 1'b0);

assign icmp_ln208_fu_758_p2 = ((add_ln207_fu_752_p2 == 32'd4) ? 1'b1 : 1'b0);

assign icmp_ln215_fu_405_p2 = ((counter_internal_blo_fu_120 < 32'd2015) ? 1'b1 : 1'b0);

assign icmp_ln224_fu_491_p2 = ((add_ln223_fu_485_p2 == 32'd8) ? 1'b1 : 1'b0);

assign icmp_ln227_fu_508_p2 = ((add_ln226_fu_502_p2 == 32'd3) ? 1'b1 : 1'b0);

assign icmp_ln230_fu_519_p2 = ((add_ln216_fu_427_p2 == 32'd3) ? 1'b1 : 1'b0);

assign icmp_ln233_fu_539_p2 = ((add_ln232_fu_533_p2 == 32'd28) ? 1'b1 : 1'b0);

assign icmp_ln236_fu_559_p2 = ((add_ln235_fu_553_p2 == 32'd28) ? 1'b1 : 1'b0);

assign icmp_ln245_1_fu_600_p2 = ((read_block_1_0_fu_108 < 32'd30) ? 1'b1 : 1'b0);

assign icmp_ln245_fu_594_p2 = ((counter_internal_blo_fu_120 < 32'd239) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_342_p2 = ((grp_fu_336_p2 == 32'd240) ? 1'b1 : 1'b0);

assign icmp_ln257_fu_639_p2 = ((add_ln256_fu_633_p2 == 32'd4) ? 1'b1 : 1'b0);

assign icmp_ln264_fu_705_p2 = ((add_ln263_fu_699_p2 == 32'd2015) ? 1'b1 : 1'b0);

assign inputBuf_0_V_address0 = zext_ln221_fu_465_p1;

assign inputBuf_1_V_address0 = zext_ln221_fu_465_p1;

assign inputBuf_2_V_address0 = zext_ln221_fu_465_p1;

assign inputBuf_3_V_address0 = zext_ln221_fu_465_p1;

assign out_V_V_TDATA = tmp_V_1_fu_788_p6;

assign select_ln208_fu_764_p3 = ((icmp_ln208_fu_758_p2[0:0] === 1'b1) ? 32'd0 : add_ln207_fu_752_p2);

assign select_ln236_1_fu_573_p3 = ((icmp_ln236_fu_559_p2[0:0] === 1'b1) ? 32'd0 : add_ln235_fu_553_p2);

assign select_ln236_fu_565_p3 = ((icmp_ln236_fu_559_p2[0:0] === 1'b1) ? 32'd0 : inp_15_0_fu_96);

assign select_ln252_1_fu_661_p3 = ((icmp_ln252_fu_342_p2[0:0] === 1'b1) ? 32'd0 : grp_fu_336_p2);

assign select_ln252_2_fu_669_p3 = ((icmp_ln252_fu_342_p2[0:0] === 1'b1) ? add_ln256_1_fu_627_p2 : trunc_ln197_fu_392_p1);

assign select_ln252_fu_653_p3 = ((icmp_ln252_fu_342_p2[0:0] === 1'b1) ? select_ln257_fu_645_p3 : current_block_write_s_fu_112);

assign select_ln257_fu_645_p3 = ((icmp_ln257_fu_639_p2[0:0] === 1'b1) ? 32'd0 : add_ln256_fu_633_p2);

assign select_ln264_fu_711_p3 = ((icmp_ln264_fu_705_p2[0:0] === 1'b1) ? 32'd0 : add_ln263_fu_699_p2);

assign shl_ln_fu_451_p3 = {{add_ln220_fu_445_p2}, {3'd0}};

assign trunc_ln197_fu_392_p1 = read_block_1_0_fu_108[4:0];

assign trunc_ln216_1_fu_433_p1 = current_block_write_s_fu_112[1:0];

assign trunc_ln216_fu_423_p1 = k_y_1_0_fu_92[1:0];

assign trunc_ln220_1_fu_441_p1 = ofm_x_1_0_fu_88[28:0];

assign trunc_ln220_fu_437_p1 = k_x_1_0_fu_100[28:0];

assign trunc_ln321_1_fu_620_p1 = current_block_write_s_fu_112[1:0];

assign trunc_ln321_fu_732_p1 = current_block_write_s_fu_112[1:0];

assign zext_ln202_fu_724_p1 = current_line_1_0_fu_116;

assign zext_ln221_fu_465_p1 = add_ln220_1_fu_459_p2;

assign zext_ln248_fu_612_p1 = current_line_1_0_fu_116;

assign zext_ln252_fu_677_p1 = select_ln252_2_fu_669_p3;

endmodule //ConvolutionInputGenerator_3_ConvolutionInputGene_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/89c3/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/6e26/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_9_0/synth/finn_design_StreamingFIFO_9_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_9:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_9,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_9_0,StreamingFIFO_9,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_9_0,StreamingFIFO_9,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_9,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_9_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [23 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 3, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [23 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 3, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_9 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/6405/hdl/verilog/StreamingFCLayer_Batch_5_Matrix_Vector_Activa.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingFCLayer_Batch_5_Matrix_Vector_Activa (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY,
        weight_V_V_TDATA,
        weight_V_V_TVALID,
        weight_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state5 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [31:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;
input  [31:0] weight_V_V_TDATA;
input   weight_V_V_TVALID;
output   weight_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;
reg weight_V_V_TREADY;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln248_fu_719_p2;
wire   [0:0] icmp_ln252_fu_734_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter2;
reg   [0:0] icmp_ln289_reg_2488;
reg   [0:0] icmp_ln289_reg_2488_pp0_iter1_reg;
reg    weight_V_V_TDATA_blk_n;
reg   [21:0] i_0_reg_547;
reg    ap_predicate_op173_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
reg    ap_block_state4_io;
reg    ap_block_pp0_stage0_11001;
wire   [21:0] i_fu_725_p2;
wire   [31:0] inElem_V_1_fu_963_p74;
wire   [6:0] trunc_ln321_fu_1113_p1;
wire   [0:0] icmp_ln271_fu_1480_p2;
reg   [0:0] icmp_ln271_reg_2443;
reg   [0:0] icmp_ln271_reg_2443_pp0_iter1_reg;
wire   [3:0] trunc_ln647_fu_1486_p1;
reg  signed [3:0] trunc_ln647_reg_2448;
reg  signed [3:0] p_Result_s_reg_2453;
reg  signed [3:0] p_Result_2_reg_2458;
reg  signed [3:0] p_Result_3_reg_2463;
reg  signed [3:0] p_Result_4_reg_2468;
reg  signed [3:0] p_Result_5_reg_2473;
reg  signed [3:0] p_Result_6_reg_2478;
reg  signed [3:0] p_Result_7_reg_2483;
wire   [0:0] icmp_ln289_fu_1566_p2;
wire  signed [7:0] mul_ln1352_5_fu_1723_p2;
reg  signed [7:0] mul_ln1352_5_reg_2492;
wire   [8:0] add_ln700_1_fu_1783_p2;
reg   [8:0] add_ln700_1_reg_2497;
wire   [8:0] add_ln700_3_fu_1789_p2;
reg   [8:0] add_ln700_3_reg_2502;
wire   [8:0] add_ln700_5_fu_1801_p2;
reg   [8:0] add_ln700_5_reg_2507;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
wire   [31:0] ap_phi_reg_pp0_iter0_act_m_val_V_reg_558;
reg   [31:0] ap_phi_reg_pp0_iter1_act_m_val_V_reg_558;
reg   [15:0] tmp_V_fu_228;
wire   [15:0] tmp_V_76_fu_1879_p2;
reg   [31:0] sf_1_fu_232;
wire   [31:0] sf_fu_1560_p2;
reg   [31:0] tmp_V_1_fu_236;
reg   [31:0] tmp_V_2_fu_240;
reg   [31:0] tmp_V_4_fu_244;
reg   [31:0] tmp_V_5_fu_248;
reg   [31:0] tmp_V_6_fu_252;
reg   [31:0] tmp_V_7_fu_256;
reg   [31:0] tmp_V_8_fu_260;
reg   [31:0] tmp_V_9_fu_264;
reg   [31:0] tmp_V_10_fu_268;
reg   [31:0] tmp_V_11_fu_272;
reg   [31:0] tmp_V_12_fu_276;
reg   [31:0] tmp_V_13_fu_280;
reg   [31:0] tmp_V_14_fu_284;
reg   [31:0] tmp_V_15_fu_288;
reg   [31:0] tmp_V_16_fu_292;
reg   [31:0] tmp_V_17_fu_296;
reg   [31:0] tmp_V_18_fu_300;
reg   [31:0] tmp_V_19_fu_304;
reg   [31:0] tmp_V_20_fu_308;
reg   [31:0] tmp_V_21_fu_312;
reg   [31:0] tmp_V_22_fu_316;
reg   [31:0] tmp_V_23_fu_320;
reg   [31:0] tmp_V_24_fu_324;
reg   [31:0] tmp_V_25_fu_328;
reg   [31:0] tmp_V_26_fu_332;
reg   [31:0] tmp_V_27_fu_336;
reg   [31:0] tmp_V_28_fu_340;
reg   [31:0] tmp_V_29_fu_344;
reg   [31:0] tmp_V_30_fu_348;
reg   [31:0] tmp_V_31_fu_352;
reg   [31:0] tmp_V_32_fu_356;
reg   [31:0] tmp_V_33_fu_360;
reg   [31:0] tmp_V_34_fu_364;
reg   [31:0] tmp_V_35_fu_368;
reg   [31:0] tmp_V_36_fu_372;
reg   [31:0] tmp_V_37_fu_376;
reg   [31:0] tmp_V_38_fu_380;
reg   [31:0] tmp_V_39_fu_384;
reg   [31:0] tmp_V_40_fu_388;
reg   [31:0] tmp_V_41_fu_392;
reg   [31:0] tmp_V_42_fu_396;
reg   [31:0] tmp_V_43_fu_400;
reg   [31:0] tmp_V_44_fu_404;
reg   [31:0] tmp_V_45_fu_408;
reg   [31:0] tmp_V_46_fu_412;
reg   [31:0] tmp_V_47_fu_416;
reg   [31:0] tmp_V_48_fu_420;
reg   [31:0] tmp_V_49_fu_424;
reg   [31:0] tmp_V_50_fu_428;
reg   [31:0] tmp_V_51_fu_432;
reg   [31:0] tmp_V_52_fu_436;
reg   [31:0] tmp_V_53_fu_440;
reg   [31:0] tmp_V_54_fu_444;
reg   [31:0] tmp_V_55_fu_448;
reg   [31:0] tmp_V_56_fu_452;
reg   [31:0] tmp_V_57_fu_456;
reg   [31:0] tmp_V_58_fu_460;
reg   [31:0] tmp_V_59_fu_464;
reg   [31:0] tmp_V_60_fu_468;
reg   [31:0] tmp_V_61_fu_472;
reg   [31:0] tmp_V_62_fu_476;
reg   [31:0] tmp_V_63_fu_480;
reg   [31:0] tmp_V_64_fu_484;
reg   [31:0] tmp_V_65_fu_488;
reg   [31:0] tmp_V_66_fu_492;
reg   [31:0] tmp_V_67_fu_496;
reg   [31:0] tmp_V_68_fu_500;
reg   [31:0] tmp_V_69_fu_504;
reg   [31:0] tmp_V_70_fu_508;
reg   [31:0] tmp_V_71_fu_512;
reg   [31:0] tmp_V_72_fu_516;
reg   [31:0] tmp_V_73_fu_520;
reg   [31:0] nf_2_fu_524;
wire   [31:0] nf_3_fu_1822_p3;
reg   [31:0] ap_sig_allocacmp_nf_2_load;
reg    ap_block_pp0_stage0_01001;
wire   [6:0] inElem_V_1_fu_963_p73;
wire  signed [3:0] trunc_ln647_1_fu_1577_p1;
wire  signed [7:0] mul_ln1352_fu_1588_p2;
wire  signed [3:0] arg_V_read_assign_1_fu_1598_p4;
wire  signed [7:0] mul_ln1352_1_fu_1615_p2;
wire  signed [3:0] arg_V_read_assign_2_fu_1625_p4;
wire  signed [7:0] mul_ln1352_2_fu_1642_p2;
wire  signed [3:0] arg_V_read_assign_3_fu_1652_p4;
wire  signed [7:0] mul_ln1352_3_fu_1669_p2;
wire  signed [3:0] arg_V_read_assign_4_fu_1679_p4;
wire  signed [7:0] mul_ln1352_4_fu_1696_p2;
wire  signed [3:0] arg_V_read_assign_5_fu_1706_p4;
wire  signed [3:0] arg_V_read_assign_6_fu_1729_p4;
wire  signed [7:0] mul_ln1352_6_fu_1746_p2;
wire  signed [3:0] arg_V_read_assign_7_fu_1756_p4;
wire  signed [7:0] mul_ln1352_7_fu_1773_p2;
wire  signed [8:0] sext_ln170_4_fu_1702_p1;
wire  signed [8:0] sext_ln170_5_fu_1752_p1;
wire  signed [8:0] sext_ln170_fu_1594_p1;
wire  signed [8:0] sext_ln170_3_fu_1675_p1;
wire  signed [8:0] sext_ln700_1_fu_1779_p1;
wire  signed [8:0] sext_ln170_1_fu_1621_p1;
wire  signed [8:0] sext_ln170_2_fu_1648_p1;
wire   [8:0] add_ln700_4_fu_1795_p2;
wire   [31:0] nf_fu_1810_p2;
wire   [0:0] icmp_ln301_fu_1816_p2;
wire  signed [15:0] sext_ln700_fu_1845_p1;
wire   [15:0] res_V_fu_1838_p3;
wire   [15:0] add_ln700_fu_1848_p2;
wire  signed [15:0] sext_ln700_2_fu_1854_p1;
wire  signed [9:0] sext_ln700_3_fu_1863_p1;
wire  signed [9:0] sext_ln700_4_fu_1866_p1;
wire   [9:0] add_ln700_6_fu_1869_p2;
wire   [15:0] add_ln700_2_fu_1857_p2;
wire  signed [15:0] sext_ln700_5_fu_1875_p1;
wire    ap_CS_fsm_state5;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

StreamingFCLayer_Batch_5_StreamingFCLayer_bkb #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 32 ),
    .din5_WIDTH( 32 ),
    .din6_WIDTH( 32 ),
    .din7_WIDTH( 32 ),
    .din8_WIDTH( 32 ),
    .din9_WIDTH( 32 ),
    .din10_WIDTH( 32 ),
    .din11_WIDTH( 32 ),
    .din12_WIDTH( 32 ),
    .din13_WIDTH( 32 ),
    .din14_WIDTH( 32 ),
    .din15_WIDTH( 32 ),
    .din16_WIDTH( 32 ),
    .din17_WIDTH( 32 ),
    .din18_WIDTH( 32 ),
    .din19_WIDTH( 32 ),
    .din20_WIDTH( 32 ),
    .din21_WIDTH( 32 ),
    .din22_WIDTH( 32 ),
    .din23_WIDTH( 32 ),
    .din24_WIDTH( 32 ),
    .din25_WIDTH( 32 ),
    .din26_WIDTH( 32 ),
    .din27_WIDTH( 32 ),
    .din28_WIDTH( 32 ),
    .din29_WIDTH( 32 ),
    .din30_WIDTH( 32 ),
    .din31_WIDTH( 32 ),
    .din32_WIDTH( 32 ),
    .din33_WIDTH( 32 ),
    .din34_WIDTH( 32 ),
    .din35_WIDTH( 32 ),
    .din36_WIDTH( 32 ),
    .din37_WIDTH( 32 ),
    .din38_WIDTH( 32 ),
    .din39_WIDTH( 32 ),
    .din40_WIDTH( 32 ),
    .din41_WIDTH( 32 ),
    .din42_WIDTH( 32 ),
    .din43_WIDTH( 32 ),
    .din44_WIDTH( 32 ),
    .din45_WIDTH( 32 ),
    .din46_WIDTH( 32 ),
    .din47_WIDTH( 32 ),
    .din48_WIDTH( 32 ),
    .din49_WIDTH( 32 ),
    .din50_WIDTH( 32 ),
    .din51_WIDTH( 32 ),
    .din52_WIDTH( 32 ),
    .din53_WIDTH( 32 ),
    .din54_WIDTH( 32 ),
    .din55_WIDTH( 32 ),
    .din56_WIDTH( 32 ),
    .din57_WIDTH( 32 ),
    .din58_WIDTH( 32 ),
    .din59_WIDTH( 32 ),
    .din60_WIDTH( 32 ),
    .din61_WIDTH( 32 ),
    .din62_WIDTH( 32 ),
    .din63_WIDTH( 32 ),
    .din64_WIDTH( 32 ),
    .din65_WIDTH( 32 ),
    .din66_WIDTH( 32 ),
    .din67_WIDTH( 32 ),
    .din68_WIDTH( 32 ),
    .din69_WIDTH( 32 ),
    .din70_WIDTH( 32 ),
    .din71_WIDTH( 32 ),
    .din72_WIDTH( 7 ),
    .dout_WIDTH( 32 ))
StreamingFCLayer_bkb_U1(
    .din0(tmp_V_1_fu_236),
    .din1(tmp_V_2_fu_240),
    .din2(tmp_V_4_fu_244),
    .din3(tmp_V_5_fu_248),
    .din4(tmp_V_6_fu_252),
    .din5(tmp_V_7_fu_256),
    .din6(tmp_V_8_fu_260),
    .din7(tmp_V_9_fu_264),
    .din8(tmp_V_10_fu_268),
    .din9(tmp_V_11_fu_272),
    .din10(tmp_V_12_fu_276),
    .din11(tmp_V_13_fu_280),
    .din12(tmp_V_14_fu_284),
    .din13(tmp_V_15_fu_288),
    .din14(tmp_V_16_fu_292),
    .din15(tmp_V_17_fu_296),
    .din16(tmp_V_18_fu_300),
    .din17(tmp_V_19_fu_304),
    .din18(tmp_V_20_fu_308),
    .din19(tmp_V_21_fu_312),
    .din20(tmp_V_22_fu_316),
    .din21(tmp_V_23_fu_320),
    .din22(tmp_V_24_fu_324),
    .din23(tmp_V_25_fu_328),
    .din24(tmp_V_26_fu_332),
    .din25(tmp_V_27_fu_336),
    .din26(tmp_V_28_fu_340),
    .din27(tmp_V_29_fu_344),
    .din28(tmp_V_30_fu_348),
    .din29(tmp_V_31_fu_352),
    .din30(tmp_V_32_fu_356),
    .din31(tmp_V_33_fu_360),
    .din32(tmp_V_34_fu_364),
    .din33(tmp_V_35_fu_368),
    .din34(tmp_V_36_fu_372),
    .din35(tmp_V_37_fu_376),
    .din36(tmp_V_38_fu_380),
    .din37(tmp_V_39_fu_384),
    .din38(tmp_V_40_fu_388),
    .din39(tmp_V_41_fu_392),
    .din40(tmp_V_42_fu_396),
    .din41(tmp_V_43_fu_400),
    .din42(tmp_V_44_fu_404),
    .din43(tmp_V_45_fu_408),
    .din44(tmp_V_46_fu_412),
    .din45(tmp_V_47_fu_416),
    .din46(tmp_V_48_fu_420),
    .din47(tmp_V_49_fu_424),
    .din48(tmp_V_50_fu_428),
    .din49(tmp_V_51_fu_432),
    .din50(tmp_V_52_fu_436),
    .din51(tmp_V_53_fu_440),
    .din52(tmp_V_54_fu_444),
    .din53(tmp_V_55_fu_448),
    .din54(tmp_V_56_fu_452),
    .din55(tmp_V_57_fu_456),
    .din56(tmp_V_58_fu_460),
    .din57(tmp_V_59_fu_464),
    .din58(tmp_V_60_fu_468),
    .din59(tmp_V_61_fu_472),
    .din60(tmp_V_62_fu_476),
    .din61(tmp_V_63_fu_480),
    .din62(tmp_V_64_fu_484),
    .din63(tmp_V_65_fu_488),
    .din64(tmp_V_66_fu_492),
    .din65(tmp_V_67_fu_496),
    .din66(tmp_V_68_fu_500),
    .din67(tmp_V_69_fu_504),
    .din68(tmp_V_70_fu_508),
    .din69(tmp_V_71_fu_512),
    .din70(tmp_V_72_fu_516),
    .din71(tmp_V_73_fu_520),
    .din72(inElem_V_1_fu_963_p73),
    .dout(inElem_V_1_fu_963_p74)
);

StreamingFCLayer_Batch_5_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U2(
    .din0(trunc_ln647_1_fu_1577_p1),
    .din1(trunc_ln647_reg_2448),
    .dout(mul_ln1352_fu_1588_p2)
);

StreamingFCLayer_Batch_5_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U3(
    .din0(arg_V_read_assign_1_fu_1598_p4),
    .din1(p_Result_s_reg_2453),
    .dout(mul_ln1352_1_fu_1615_p2)
);

StreamingFCLayer_Batch_5_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U4(
    .din0(arg_V_read_assign_2_fu_1625_p4),
    .din1(p_Result_2_reg_2458),
    .dout(mul_ln1352_2_fu_1642_p2)
);

StreamingFCLayer_Batch_5_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U5(
    .din0(arg_V_read_assign_3_fu_1652_p4),
    .din1(p_Result_3_reg_2463),
    .dout(mul_ln1352_3_fu_1669_p2)
);

StreamingFCLayer_Batch_5_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U6(
    .din0(arg_V_read_assign_4_fu_1679_p4),
    .din1(p_Result_4_reg_2468),
    .dout(mul_ln1352_4_fu_1696_p2)
);

StreamingFCLayer_Batch_5_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U7(
    .din0(arg_V_read_assign_5_fu_1706_p4),
    .din1(p_Result_5_reg_2473),
    .dout(mul_ln1352_5_fu_1723_p2)
);

StreamingFCLayer_Batch_5_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U8(
    .din0(arg_V_read_assign_6_fu_1729_p4),
    .din1(p_Result_6_reg_2478),
    .dout(mul_ln1352_6_fu_1746_p2)
);

StreamingFCLayer_Batch_5_StreamingFCLayer_cud #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_cud_U9(
    .din0(arg_V_read_assign_7_fu_1756_p4),
    .din1(p_Result_7_reg_2483),
    .dout(mul_ln1352_7_fu_1773_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd0) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_558 <= inElem_V_1_fu_963_p74;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd70)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd69)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd68)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd67)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd66)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd65)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd64)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd63)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd62)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd61)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd60)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd59)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd58)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd57)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd56)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd55)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd54)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd53)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd52)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd51)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd50)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd49)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd48)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd47)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd46)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd45)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd44)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd43)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd42)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd41)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd40)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd39)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd38)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd37)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd36)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd35)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd34)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd33)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd32)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd31)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd30)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd29)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd28)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd27)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd26)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd25)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd24)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd23)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd22)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd21)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd20)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd19)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd18)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd17)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd16)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd15)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd14)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd13)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd12)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd11)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd10)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd9)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd8)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd7)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd6)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd5)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd4)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd3)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd2)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd1)) | (~(trunc_ln321_fu_1113_p1 == 7'd70) & ~(trunc_ln321_fu_1113_p1 == 7'd69) & ~(trunc_ln321_fu_1113_p1 == 7'd68) & ~(trunc_ln321_fu_1113_p1 == 7'd67) & ~(trunc_ln321_fu_1113_p1 == 7'd66) & ~(trunc_ln321_fu_1113_p1 == 7'd65) & ~(trunc_ln321_fu_1113_p1 == 7'd64) & ~(trunc_ln321_fu_1113_p1 == 7'd63) & ~(trunc_ln321_fu_1113_p1 == 7'd62) & ~(trunc_ln321_fu_1113_p1 == 7'd61) & ~(trunc_ln321_fu_1113_p1 == 7'd60) & ~(trunc_ln321_fu_1113_p1 == 7'd59) & ~(trunc_ln321_fu_1113_p1 == 7'd58) & ~(trunc_ln321_fu_1113_p1 == 7'd57) & ~(trunc_ln321_fu_1113_p1 == 7'd56) & ~(trunc_ln321_fu_1113_p1 == 7'd55) & ~(trunc_ln321_fu_1113_p1 == 7'd54) & ~(trunc_ln321_fu_1113_p1 == 7'd53) & ~(trunc_ln321_fu_1113_p1 == 7'd52) & ~(trunc_ln321_fu_1113_p1 == 7'd51) & ~(trunc_ln321_fu_1113_p1 == 7'd50) & ~(trunc_ln321_fu_1113_p1 == 7'd49) & ~(trunc_ln321_fu_1113_p1 == 7'd48) & ~(trunc_ln321_fu_1113_p1 == 7'd47) & ~(trunc_ln321_fu_1113_p1 == 7'd46) & ~(trunc_ln321_fu_1113_p1 == 7'd45) & ~(trunc_ln321_fu_1113_p1 == 7'd44) & ~(trunc_ln321_fu_1113_p1 == 7'd43) & ~(trunc_ln321_fu_1113_p1 == 7'd42) & ~(trunc_ln321_fu_1113_p1 == 7'd41) & ~(trunc_ln321_fu_1113_p1 == 7'd40) & ~(trunc_ln321_fu_1113_p1 == 7'd39) & ~(trunc_ln321_fu_1113_p1 == 7'd38) & ~(trunc_ln321_fu_1113_p1 == 7'd37) & ~(trunc_ln321_fu_1113_p1 == 7'd36) & ~(trunc_ln321_fu_1113_p1 == 7'd35) & ~(trunc_ln321_fu_1113_p1 == 7'd34) & ~(trunc_ln321_fu_1113_p1 == 7'd33) & ~(trunc_ln321_fu_1113_p1 == 7'd32) & ~(trunc_ln321_fu_1113_p1 == 7'd31) & ~(trunc_ln321_fu_1113_p1 == 7'd30) & ~(trunc_ln321_fu_1113_p1 == 7'd29) & ~(trunc_ln321_fu_1113_p1 == 7'd28) & ~(trunc_ln321_fu_1113_p1 == 7'd27) & ~(trunc_ln321_fu_1113_p1 == 7'd26) & ~(trunc_ln321_fu_1113_p1 == 7'd25) & ~(trunc_ln321_fu_1113_p1 == 7'd24) & ~(trunc_ln321_fu_1113_p1 == 7'd23) & ~(trunc_ln321_fu_1113_p1 == 7'd22) & ~(trunc_ln321_fu_1113_p1 == 7'd21) & ~(trunc_ln321_fu_1113_p1 == 7'd20) & ~(trunc_ln321_fu_1113_p1 == 7'd19) & ~(trunc_ln321_fu_1113_p1 == 7'd18) & ~(trunc_ln321_fu_1113_p1 == 7'd17) & ~(trunc_ln321_fu_1113_p1 == 7'd16) & ~(trunc_ln321_fu_1113_p1 == 7'd15) & ~(trunc_ln321_fu_1113_p1 == 7'd14) & ~(trunc_ln321_fu_1113_p1 == 7'd13) & ~(trunc_ln321_fu_1113_p1 == 7'd12) & ~(trunc_ln321_fu_1113_p1 == 7'd11) & ~(trunc_ln321_fu_1113_p1 == 7'd10) & ~(trunc_ln321_fu_1113_p1 == 7'd9) & ~(trunc_ln321_fu_1113_p1 == 7'd8) & ~(trunc_ln321_fu_1113_p1 == 7'd7) & ~(trunc_ln321_fu_1113_p1 == 7'd6) & ~(trunc_ln321_fu_1113_p1 == 7'd5) & ~(trunc_ln321_fu_1113_p1 == 7'd4) & ~(trunc_ln321_fu_1113_p1 == 7'd3) & ~(trunc_ln321_fu_1113_p1 == 7'd2) & ~(trunc_ln321_fu_1113_p1 == 7'd1) & ~(trunc_ln321_fu_1113_p1 == 7'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd0)))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_558 <= in_V_V_TDATA;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_558 <= ap_phi_reg_pp0_iter0_act_m_val_V_reg_558;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_reg_547 <= i_fu_725_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_reg_547 <= 22'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_2488 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        nf_2_fu_524 <= nf_3_fu_1822_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        nf_2_fu_524 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_1566_p2 == 1'd0) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        sf_1_fu_232 <= sf_fu_1560_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_1566_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        sf_1_fu_232 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln700_1_reg_2497 <= add_ln700_1_fu_1783_p2;
        add_ln700_3_reg_2502 <= add_ln700_3_fu_1789_p2;
        add_ln700_5_reg_2507 <= add_ln700_5_fu_1801_p2;
        icmp_ln271_reg_2443_pp0_iter1_reg <= icmp_ln271_reg_2443;
        icmp_ln289_reg_2488_pp0_iter1_reg <= icmp_ln289_reg_2488;
        mul_ln1352_5_reg_2492 <= mul_ln1352_5_fu_1723_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_719_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln271_reg_2443 <= icmp_ln271_fu_1480_p2;
        icmp_ln289_reg_2488 <= icmp_ln289_fu_1566_p2;
        p_Result_2_reg_2458 <= {{weight_V_V_TDATA[11:8]}};
        p_Result_3_reg_2463 <= {{weight_V_V_TDATA[15:12]}};
        p_Result_4_reg_2468 <= {{weight_V_V_TDATA[19:16]}};
        p_Result_5_reg_2473 <= {{weight_V_V_TDATA[23:20]}};
        p_Result_6_reg_2478 <= {{weight_V_V_TDATA[27:24]}};
        p_Result_7_reg_2483 <= {{weight_V_V_TDATA[31:28]}};
        p_Result_s_reg_2453 <= {{weight_V_V_TDATA[7:4]}};
        trunc_ln647_reg_2448 <= trunc_ln647_fu_1486_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd8))) begin
        tmp_V_10_fu_268 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd9))) begin
        tmp_V_11_fu_272 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd10))) begin
        tmp_V_12_fu_276 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd11))) begin
        tmp_V_13_fu_280 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd12))) begin
        tmp_V_14_fu_284 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd13))) begin
        tmp_V_15_fu_288 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd14))) begin
        tmp_V_16_fu_292 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd15))) begin
        tmp_V_17_fu_296 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd16))) begin
        tmp_V_18_fu_300 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd17))) begin
        tmp_V_19_fu_304 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd0))) begin
        tmp_V_1_fu_236 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd18))) begin
        tmp_V_20_fu_308 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd19))) begin
        tmp_V_21_fu_312 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd20))) begin
        tmp_V_22_fu_316 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd21))) begin
        tmp_V_23_fu_320 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd22))) begin
        tmp_V_24_fu_324 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd23))) begin
        tmp_V_25_fu_328 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd24))) begin
        tmp_V_26_fu_332 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd25))) begin
        tmp_V_27_fu_336 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd26))) begin
        tmp_V_28_fu_340 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd27))) begin
        tmp_V_29_fu_344 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd1))) begin
        tmp_V_2_fu_240 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd28))) begin
        tmp_V_30_fu_348 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd29))) begin
        tmp_V_31_fu_352 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd30))) begin
        tmp_V_32_fu_356 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd31))) begin
        tmp_V_33_fu_360 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd32))) begin
        tmp_V_34_fu_364 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd33))) begin
        tmp_V_35_fu_368 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd34))) begin
        tmp_V_36_fu_372 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd35))) begin
        tmp_V_37_fu_376 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd36))) begin
        tmp_V_38_fu_380 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd37))) begin
        tmp_V_39_fu_384 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd38))) begin
        tmp_V_40_fu_388 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd39))) begin
        tmp_V_41_fu_392 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd40))) begin
        tmp_V_42_fu_396 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd41))) begin
        tmp_V_43_fu_400 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd42))) begin
        tmp_V_44_fu_404 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd43))) begin
        tmp_V_45_fu_408 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd44))) begin
        tmp_V_46_fu_412 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd45))) begin
        tmp_V_47_fu_416 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd46))) begin
        tmp_V_48_fu_420 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd47))) begin
        tmp_V_49_fu_424 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd2))) begin
        tmp_V_4_fu_244 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd48))) begin
        tmp_V_50_fu_428 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd49))) begin
        tmp_V_51_fu_432 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd50))) begin
        tmp_V_52_fu_436 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd51))) begin
        tmp_V_53_fu_440 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd52))) begin
        tmp_V_54_fu_444 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd53))) begin
        tmp_V_55_fu_448 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd54))) begin
        tmp_V_56_fu_452 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd55))) begin
        tmp_V_57_fu_456 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd56))) begin
        tmp_V_58_fu_460 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd57))) begin
        tmp_V_59_fu_464 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd3))) begin
        tmp_V_5_fu_248 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd58))) begin
        tmp_V_60_fu_468 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd59))) begin
        tmp_V_61_fu_472 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd60))) begin
        tmp_V_62_fu_476 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd61))) begin
        tmp_V_63_fu_480 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd62))) begin
        tmp_V_64_fu_484 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd63))) begin
        tmp_V_65_fu_488 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd64))) begin
        tmp_V_66_fu_492 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd65))) begin
        tmp_V_67_fu_496 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd66))) begin
        tmp_V_68_fu_500 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd67))) begin
        tmp_V_69_fu_504 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd4))) begin
        tmp_V_6_fu_252 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd68))) begin
        tmp_V_70_fu_508 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd69))) begin
        tmp_V_71_fu_512 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd70))) begin
        tmp_V_72_fu_516 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if ((~(trunc_ln321_fu_1113_p1 == 7'd70) & ~(trunc_ln321_fu_1113_p1 == 7'd69) & ~(trunc_ln321_fu_1113_p1 == 7'd68) & ~(trunc_ln321_fu_1113_p1 == 7'd67) & ~(trunc_ln321_fu_1113_p1 == 7'd66) & ~(trunc_ln321_fu_1113_p1 == 7'd65) & ~(trunc_ln321_fu_1113_p1 == 7'd64) & ~(trunc_ln321_fu_1113_p1 == 7'd63) & ~(trunc_ln321_fu_1113_p1 == 7'd62) & ~(trunc_ln321_fu_1113_p1 == 7'd61) & ~(trunc_ln321_fu_1113_p1 == 7'd60) & ~(trunc_ln321_fu_1113_p1 == 7'd59) & ~(trunc_ln321_fu_1113_p1 == 7'd58) & ~(trunc_ln321_fu_1113_p1 == 7'd57) & ~(trunc_ln321_fu_1113_p1 == 7'd56) & ~(trunc_ln321_fu_1113_p1 == 7'd55) & ~(trunc_ln321_fu_1113_p1 == 7'd54) & ~(trunc_ln321_fu_1113_p1 == 7'd53) & ~(trunc_ln321_fu_1113_p1 == 7'd52) & ~(trunc_ln321_fu_1113_p1 == 7'd51) & ~(trunc_ln321_fu_1113_p1 == 7'd50) & ~(trunc_ln321_fu_1113_p1 == 7'd49) & ~(trunc_ln321_fu_1113_p1 == 7'd48) & ~(trunc_ln321_fu_1113_p1 == 7'd47) & ~(trunc_ln321_fu_1113_p1 == 7'd46) & ~(trunc_ln321_fu_1113_p1 == 7'd45) & ~(trunc_ln321_fu_1113_p1 == 7'd44) & ~(trunc_ln321_fu_1113_p1 == 7'd43) & ~(trunc_ln321_fu_1113_p1 == 7'd42) & ~(trunc_ln321_fu_1113_p1 == 7'd41) & ~(trunc_ln321_fu_1113_p1 == 7'd40) & ~(trunc_ln321_fu_1113_p1 == 7'd39) & ~(trunc_ln321_fu_1113_p1 == 7'd38) & ~(trunc_ln321_fu_1113_p1 == 7'd37) & ~(trunc_ln321_fu_1113_p1 == 7'd36) & ~(trunc_ln321_fu_1113_p1 == 7'd35) & ~(trunc_ln321_fu_1113_p1 == 7'd34) & ~(trunc_ln321_fu_1113_p1 == 7'd33) & ~(trunc_ln321_fu_1113_p1 == 7'd32) & ~(trunc_ln321_fu_1113_p1 == 7'd31) & ~(trunc_ln321_fu_1113_p1 == 7'd30) & ~(trunc_ln321_fu_1113_p1 == 7'd29) & ~(trunc_ln321_fu_1113_p1 == 7'd28) & ~(trunc_ln321_fu_1113_p1 == 7'd27) & ~(trunc_ln321_fu_1113_p1 == 7'd26) & ~(trunc_ln321_fu_1113_p1 == 7'd25) & ~(trunc_ln321_fu_1113_p1 == 7'd24) & ~(trunc_ln321_fu_1113_p1 == 7'd23) & ~(trunc_ln321_fu_1113_p1 == 7'd22) & ~(trunc_ln321_fu_1113_p1 == 7'd21) & ~(trunc_ln321_fu_1113_p1 == 7'd20) & ~(trunc_ln321_fu_1113_p1 == 7'd19) & ~(trunc_ln321_fu_1113_p1 == 7'd18) & ~(trunc_ln321_fu_1113_p1 == 7'd17) & ~(trunc_ln321_fu_1113_p1 == 7'd16) & ~(trunc_ln321_fu_1113_p1 == 7'd15) & ~(trunc_ln321_fu_1113_p1 == 7'd14) & ~(trunc_ln321_fu_1113_p1 == 7'd13) & ~(trunc_ln321_fu_1113_p1 == 7'd12) & ~(trunc_ln321_fu_1113_p1 == 7'd11) & ~(trunc_ln321_fu_1113_p1 == 7'd10) & ~(trunc_ln321_fu_1113_p1 == 7'd9) & ~(trunc_ln321_fu_1113_p1 == 7'd8) & ~(trunc_ln321_fu_1113_p1 == 7'd7) & ~(trunc_ln321_fu_1113_p1 == 7'd6) & ~(trunc_ln321_fu_1113_p1 == 7'd5) & ~(trunc_ln321_fu_1113_p1 == 7'd4) & ~(trunc_ln321_fu_1113_p1 == 7'd3) & ~(trunc_ln321_fu_1113_p1 == 7'd2) & ~(trunc_ln321_fu_1113_p1 == 7'd1) & ~(trunc_ln321_fu_1113_p1 == 7'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_73_fu_520 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd5))) begin
        tmp_V_7_fu_256 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd6))) begin
        tmp_V_8_fu_260 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (trunc_ln321_fu_1113_p1 == 7'd7))) begin
        tmp_V_9_fu_264 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        tmp_V_fu_228 <= tmp_V_76_fu_1879_p2;
    end
end

always @ (*) begin
    if ((icmp_ln248_fu_719_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state5) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state5)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_2488 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_sig_allocacmp_nf_2_load = nf_3_fu_1822_p3;
    end else begin
        ap_sig_allocacmp_nf_2_load = nf_2_fu_524;
    end
end

always @ (*) begin
    if (((icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op173_read_state2 == 1'b1))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_2488_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_2488_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln248_fu_719_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TDATA_blk_n = weight_V_V_TVALID;
    end else begin
        weight_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_719_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TREADY = 1'b1;
    end else begin
        weight_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln248_fu_719_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)) & ~((ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)) | ((icmp_ln248_fu_719_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln700_1_fu_1783_p2 = ($signed(sext_ln170_4_fu_1702_p1) + $signed(sext_ln170_5_fu_1752_p1));

assign add_ln700_2_fu_1857_p2 = ($signed(add_ln700_fu_1848_p2) + $signed(sext_ln700_2_fu_1854_p1));

assign add_ln700_3_fu_1789_p2 = ($signed(sext_ln170_fu_1594_p1) + $signed(sext_ln170_3_fu_1675_p1));

assign add_ln700_4_fu_1795_p2 = ($signed(sext_ln700_1_fu_1779_p1) + $signed(sext_ln170_1_fu_1621_p1));

assign add_ln700_5_fu_1801_p2 = ($signed(sext_ln170_2_fu_1648_p1) + $signed(add_ln700_4_fu_1795_p2));

assign add_ln700_6_fu_1869_p2 = ($signed(sext_ln700_3_fu_1863_p1) + $signed(sext_ln700_4_fu_1866_p1));

assign add_ln700_fu_1848_p2 = ($signed(sext_ln700_fu_1845_p1) + $signed(res_V_fu_1838_p3));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state5 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op173_read_state2 == 1'b1)) | ((icmp_ln248_fu_719_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_block_state4_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op173_read_state2 == 1'b1)) | ((icmp_ln248_fu_719_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_block_state4_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op173_read_state2 == 1'b1)) | ((icmp_ln248_fu_719_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op173_read_state2 == 1'b1)) | ((icmp_ln248_fu_719_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state4_io = ((icmp_ln289_reg_2488_pp0_iter1_reg == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_reg_pp0_iter0_act_m_val_V_reg_558 = 'bx;

always @ (*) begin
    ap_predicate_op173_read_state2 = ((icmp_ln252_fu_734_p2 == 1'd1) & (icmp_ln248_fu_719_p2 == 1'd0));
end

assign arg_V_read_assign_1_fu_1598_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_558[7:4]}};

assign arg_V_read_assign_2_fu_1625_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_558[11:8]}};

assign arg_V_read_assign_3_fu_1652_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_558[15:12]}};

assign arg_V_read_assign_4_fu_1679_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_558[19:16]}};

assign arg_V_read_assign_5_fu_1706_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_558[23:20]}};

assign arg_V_read_assign_6_fu_1729_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_558[27:24]}};

assign arg_V_read_assign_7_fu_1756_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_558[31:28]}};

assign i_fu_725_p2 = (i_0_reg_547 + 22'd1);

assign icmp_ln248_fu_719_p2 = ((i_0_reg_547 == 22'd3612672) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_734_p2 = ((ap_sig_allocacmp_nf_2_load == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln271_fu_1480_p2 = ((sf_1_fu_232 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln289_fu_1566_p2 = ((sf_fu_1560_p2 == 32'd72) ? 1'b1 : 1'b0);

assign icmp_ln301_fu_1816_p2 = ((nf_fu_1810_p2 == 32'd64) ? 1'b1 : 1'b0);

assign inElem_V_1_fu_963_p73 = sf_1_fu_232[6:0];

assign nf_3_fu_1822_p3 = ((icmp_ln301_fu_1816_p2[0:0] === 1'b1) ? 32'd0 : nf_fu_1810_p2);

assign nf_fu_1810_p2 = (nf_2_fu_524 + 32'd1);

assign out_V_V_TDATA = ($signed(add_ln700_2_fu_1857_p2) + $signed(sext_ln700_5_fu_1875_p1));

assign res_V_fu_1838_p3 = ((icmp_ln271_reg_2443_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : tmp_V_fu_228);

assign sext_ln170_1_fu_1621_p1 = mul_ln1352_1_fu_1615_p2;

assign sext_ln170_2_fu_1648_p1 = mul_ln1352_2_fu_1642_p2;

assign sext_ln170_3_fu_1675_p1 = mul_ln1352_3_fu_1669_p2;

assign sext_ln170_4_fu_1702_p1 = mul_ln1352_4_fu_1696_p2;

assign sext_ln170_5_fu_1752_p1 = mul_ln1352_6_fu_1746_p2;

assign sext_ln170_fu_1594_p1 = mul_ln1352_fu_1588_p2;

assign sext_ln700_1_fu_1779_p1 = mul_ln1352_7_fu_1773_p2;

assign sext_ln700_2_fu_1854_p1 = $signed(add_ln700_1_reg_2497);

assign sext_ln700_3_fu_1863_p1 = $signed(add_ln700_3_reg_2502);

assign sext_ln700_4_fu_1866_p1 = $signed(add_ln700_5_reg_2507);

assign sext_ln700_5_fu_1875_p1 = $signed(add_ln700_6_fu_1869_p2);

assign sext_ln700_fu_1845_p1 = mul_ln1352_5_reg_2492;

assign sf_fu_1560_p2 = (32'd1 + sf_1_fu_232);

assign tmp_V_76_fu_1879_p2 = ($signed(add_ln700_2_fu_1857_p2) + $signed(sext_ln700_5_fu_1875_p1));

assign trunc_ln321_fu_1113_p1 = sf_1_fu_232[6:0];

assign trunc_ln647_1_fu_1577_p1 = ap_phi_reg_pp0_iter1_act_m_val_V_reg_558[3:0];

assign trunc_ln647_fu_1486_p1 = weight_V_V_TDATA[3:0];

endmodule //StreamingFCLayer_Batch_5_Matrix_Vector_Activa
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/db73/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc0C.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcc0C_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc0C_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcc0C(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcc0C_rom Thresholding_Batch_0_Thresholding_Batcc0C_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActShg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActShg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActShg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActShg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActShg_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActShg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcqcK.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcqcK_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 5;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcqcK_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcqcK(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd5;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcqcK_rom Thresholding_Batch_0_Thresholding_BatcqcK_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbll.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbll_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbll_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbll(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbll_rom Thresholding_Batch_0_Thresholding_Batcbll_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActpcA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActpcA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActpcA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActpcA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActpcA_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActpcA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/a3f1/hdl/verilog/ConvolutionInputGenerator_1_ConvolutionInputGene_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module ConvolutionInputGenerator_1_ConvolutionInputGene_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [15:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln197_fu_368_p2;
wire   [0:0] icmp_ln199_fu_390_p2;
wire   [0:0] and_ln245_fu_600_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln199_reg_887;
reg   [0:0] icmp_ln215_reg_891;
reg   [10:0] i_0_0_reg_271;
reg    ap_predicate_op119_read_state2;
reg    ap_predicate_op162_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_predicate_op205_write_state3;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [10:0] add_ln197_fu_374_p2;
wire   [0:0] icmp_ln215_fu_399_p2;
wire   [1:0] add_ln221_fu_473_p2;
reg   [1:0] add_ln221_reg_895;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
wire   [7:0] inputBuf_0_V_address0;
reg    inputBuf_0_V_ce0;
wire   [15:0] inputBuf_0_V_q0;
reg   [7:0] inputBuf_0_V_address1;
reg    inputBuf_0_V_ce1;
reg    inputBuf_0_V_we1;
wire   [7:0] inputBuf_1_V_address0;
reg    inputBuf_1_V_ce0;
wire   [15:0] inputBuf_1_V_q0;
reg   [7:0] inputBuf_1_V_address1;
reg    inputBuf_1_V_ce1;
reg    inputBuf_1_V_we1;
wire   [7:0] inputBuf_2_V_address0;
reg    inputBuf_2_V_ce0;
wire   [15:0] inputBuf_2_V_q0;
reg   [7:0] inputBuf_2_V_address1;
reg    inputBuf_2_V_ce1;
reg    inputBuf_2_V_we1;
wire   [7:0] inputBuf_3_V_address0;
reg    inputBuf_3_V_ce0;
wire   [15:0] inputBuf_3_V_q0;
reg   [7:0] inputBuf_3_V_address1;
reg    inputBuf_3_V_ce1;
reg    inputBuf_3_V_we1;
wire   [63:0] zext_ln221_fu_459_p1;
wire   [63:0] zext_ln248_fu_606_p1;
wire   [63:0] zext_ln202_fu_718_p1;
reg   [31:0] ofm_y_1_0_fu_78;
wire   [31:0] select_ln236_1_fu_567_p3;
wire   [0:0] icmp_ln224_fu_485_p2;
wire   [0:0] icmp_ln227_fu_502_p2;
wire   [0:0] icmp_ln230_fu_513_p2;
wire   [0:0] icmp_ln233_fu_533_p2;
reg   [31:0] ofm_x_1_0_fu_82;
wire   [31:0] add_ln232_fu_527_p2;
reg   [31:0] k_y_1_0_fu_86;
wire   [31:0] add_ln216_fu_421_p2;
reg   [31:0] inp_15_0_fu_90;
wire   [31:0] select_ln236_fu_559_p3;
wire   [31:0] add_ln204_fu_730_p2;
reg   [31:0] k_x_1_0_fu_94;
wire   [31:0] add_ln226_fu_496_p2;
reg   [31:0] count_simd_1_0_fu_98;
wire   [31:0] add_ln223_fu_479_p2;
reg   [31:0] read_block_1_0_fu_102;
wire   [31:0] zext_ln252_fu_671_p1;
wire   [31:0] add_ln211_fu_766_p2;
wire   [0:0] icmp_ln205_fu_342_p2;
reg   [31:0] current_block_write_s_fu_106;
wire   [31:0] select_ln252_fu_647_p3;
wire   [31:0] select_ln208_fu_758_p3;
reg   [31:0] current_line_1_0_fu_110;
wire   [31:0] select_ln252_1_fu_655_p3;
wire   [31:0] grp_fu_330_p2;
reg   [31:0] counter_internal_blo_fu_114;
wire   [31:0] select_ln264_fu_705_p3;
wire   [15:0] tmp_V_1_fu_782_p6;
reg    ap_block_pp0_stage0_01001;
wire   [1:0] trunc_ln321_1_fu_614_p1;
wire   [1:0] trunc_ln321_fu_726_p1;
wire   [25:0] trunc_ln220_1_fu_435_p1;
wire   [25:0] trunc_ln220_fu_431_p1;
wire   [25:0] add_ln220_fu_439_p2;
wire   [31:0] shl_ln_fu_445_p3;
wire   [31:0] add_ln220_1_fu_453_p2;
wire   [1:0] trunc_ln216_1_fu_427_p1;
wire   [1:0] add_ln221_1_fu_467_p2;
wire   [1:0] trunc_ln216_fu_417_p1;
wire   [0:0] icmp_ln236_fu_553_p2;
wire   [31:0] add_ln235_fu_547_p2;
wire   [0:0] icmp_ln245_fu_588_p2;
wire   [0:0] icmp_ln245_1_fu_594_p2;
wire   [1:0] trunc_ln197_fu_386_p1;
wire   [31:0] add_ln256_fu_627_p2;
wire   [0:0] icmp_ln257_fu_633_p2;
wire   [0:0] icmp_ln252_fu_336_p2;
wire   [31:0] select_ln257_fu_639_p3;
wire   [1:0] add_ln256_1_fu_621_p2;
wire   [1:0] select_ln252_2_fu_663_p3;
wire   [31:0] add_ln263_fu_693_p2;
wire   [0:0] icmp_ln264_fu_699_p2;
wire   [31:0] add_ln207_fu_746_p2;
wire   [0:0] icmp_ln208_fu_752_p2;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_block_pp0;
reg    ap_predicate_op127_store_state2;
reg    ap_enable_operation_127;
reg    ap_enable_state2_pp0_iter0_stage0;
reg    ap_predicate_op69_load_state2;
reg    ap_enable_operation_69;
reg    ap_predicate_op202_load_state3;
reg    ap_enable_operation_202;
reg    ap_enable_state3_pp0_iter1_stage0;
reg    ap_predicate_op170_store_state2;
reg    ap_enable_operation_170;
reg    ap_predicate_op129_store_state2;
reg    ap_enable_operation_129;
reg    ap_predicate_op67_load_state2;
reg    ap_enable_operation_67;
reg    ap_predicate_op201_load_state3;
reg    ap_enable_operation_201;
reg    ap_predicate_op172_store_state2;
reg    ap_enable_operation_172;
reg    ap_predicate_op131_store_state2;
reg    ap_enable_operation_131;
reg    ap_predicate_op65_load_state2;
reg    ap_enable_operation_65;
reg    ap_predicate_op200_load_state3;
reg    ap_enable_operation_200;
reg    ap_predicate_op174_store_state2;
reg    ap_enable_operation_174;
reg    ap_predicate_op133_store_state2;
reg    ap_enable_operation_133;
reg    ap_predicate_op71_load_state2;
reg    ap_enable_operation_71;
reg    ap_predicate_op203_load_state3;
reg    ap_enable_operation_203;
reg    ap_predicate_op176_store_state2;
reg    ap_enable_operation_176;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_657;
reg    ap_condition_230;
reg    ap_condition_663;
reg    ap_condition_667;
reg    ap_condition_671;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

ConvolutionInputGenerator_1_ConvolutionInputGbkb #(
    .DataWidth( 16 ),
    .AddressRange( 192 ),
    .AddressWidth( 8 ))
inputBuf_0_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_0_V_address0),
    .ce0(inputBuf_0_V_ce0),
    .q0(inputBuf_0_V_q0),
    .address1(inputBuf_0_V_address1),
    .ce1(inputBuf_0_V_ce1),
    .we1(inputBuf_0_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_1_ConvolutionInputGbkb #(
    .DataWidth( 16 ),
    .AddressRange( 192 ),
    .AddressWidth( 8 ))
inputBuf_1_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_1_V_address0),
    .ce0(inputBuf_1_V_ce0),
    .q0(inputBuf_1_V_q0),
    .address1(inputBuf_1_V_address1),
    .ce1(inputBuf_1_V_ce1),
    .we1(inputBuf_1_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_1_ConvolutionInputGbkb #(
    .DataWidth( 16 ),
    .AddressRange( 192 ),
    .AddressWidth( 8 ))
inputBuf_2_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_2_V_address0),
    .ce0(inputBuf_2_V_ce0),
    .q0(inputBuf_2_V_q0),
    .address1(inputBuf_2_V_address1),
    .ce1(inputBuf_2_V_ce1),
    .we1(inputBuf_2_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_1_ConvolutionInputGbkb #(
    .DataWidth( 16 ),
    .AddressRange( 192 ),
    .AddressWidth( 8 ))
inputBuf_3_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_3_V_address0),
    .ce0(inputBuf_3_V_ce0),
    .q0(inputBuf_3_V_q0),
    .address1(inputBuf_3_V_address1),
    .ce1(inputBuf_3_V_ce1),
    .we1(inputBuf_3_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_1_ConvolutionInputGfYi #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .din2_WIDTH( 16 ),
    .din3_WIDTH( 16 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 16 ))
ConvolutionInputGfYi_U1(
    .din0(inputBuf_0_V_q0),
    .din1(inputBuf_1_V_q0),
    .din2(inputBuf_2_V_q0),
    .din3(inputBuf_3_V_q0),
    .din4(add_ln221_reg_895),
    .dout(tmp_V_1_fu_782_p6)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln224_fu_485_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        count_simd_1_0_fu_98 <= add_ln223_fu_479_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln227_fu_502_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln230_fu_513_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln230_fu_513_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln233_fu_533_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln233_fu_533_p2 == 1'd1) & (icmp_ln230_fu_513_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        count_simd_1_0_fu_98 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        counter_internal_blo_fu_114 <= select_ln264_fu_705_p3;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_342_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        counter_internal_blo_fu_114 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_342_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_block_write_s_fu_106 <= select_ln208_fu_758_p3;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_block_write_s_fu_106 <= select_ln252_fu_647_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        current_block_write_s_fu_106 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln205_fu_342_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_line_1_0_fu_110 <= grp_fu_330_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_line_1_0_fu_110 <= select_ln252_1_fu_655_p3;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_342_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        current_line_1_0_fu_110 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_0_reg_271 <= 11'd0;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_0_reg_271 <= add_ln197_fu_374_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inp_15_0_fu_90 <= add_ln204_fu_730_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln233_fu_533_p2 == 1'd1) & (icmp_ln230_fu_513_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inp_15_0_fu_90 <= select_ln236_fu_559_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        inp_15_0_fu_90 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln227_fu_502_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        k_x_1_0_fu_94 <= add_ln226_fu_496_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln230_fu_513_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln230_fu_513_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln233_fu_533_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln233_fu_533_p2 == 1'd1) & (icmp_ln230_fu_513_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        k_x_1_0_fu_94 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln230_fu_513_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        k_y_1_0_fu_86 <= add_ln216_fu_421_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln230_fu_513_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        k_y_1_0_fu_86 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln230_fu_513_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln233_fu_533_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ofm_x_1_0_fu_82 <= add_ln232_fu_527_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln233_fu_533_p2 == 1'd1) & (icmp_ln230_fu_513_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ofm_x_1_0_fu_82 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln233_fu_533_p2 == 1'd1) & (icmp_ln230_fu_513_p2 == 1'd1) & (icmp_ln227_fu_502_p2 == 1'd1) & (icmp_ln224_fu_485_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ofm_y_1_0_fu_78 <= select_ln236_1_fu_567_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        ofm_y_1_0_fu_78 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_342_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        read_block_1_0_fu_102 <= add_ln211_fu_766_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        read_block_1_0_fu_102 <= zext_ln252_fu_671_p1;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        read_block_1_0_fu_102 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln221_reg_895 <= add_ln221_fu_473_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln197_fu_368_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln199_reg_887 <= icmp_ln199_fu_390_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln215_reg_891 <= icmp_ln215_fu_399_p2;
    end
end

always @ (*) begin
    if ((icmp_ln197_fu_368_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op119_read_state2 == 1'b1)))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_390_p2 == 1'd1) & (trunc_ln321_fu_726_p1 == 2'd0))) begin
            inputBuf_0_V_address1 = zext_ln202_fu_718_p1;
        end else if ((1'b1 == ap_condition_657)) begin
            inputBuf_0_V_address1 = zext_ln248_fu_606_p1;
        end else begin
            inputBuf_0_V_address1 = 'bx;
        end
    end else begin
        inputBuf_0_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_0_V_ce0 = 1'b1;
    end else begin
        inputBuf_0_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_0_V_ce1 = 1'b1;
    end else begin
        inputBuf_0_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_0_V_we1 = 1'b1;
    end else begin
        inputBuf_0_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_390_p2 == 1'd1) & (trunc_ln321_fu_726_p1 == 2'd1))) begin
            inputBuf_1_V_address1 = zext_ln202_fu_718_p1;
        end else if ((1'b1 == ap_condition_663)) begin
            inputBuf_1_V_address1 = zext_ln248_fu_606_p1;
        end else begin
            inputBuf_1_V_address1 = 'bx;
        end
    end else begin
        inputBuf_1_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_1_V_ce0 = 1'b1;
    end else begin
        inputBuf_1_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_1_V_ce1 = 1'b1;
    end else begin
        inputBuf_1_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_1_V_we1 = 1'b1;
    end else begin
        inputBuf_1_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_390_p2 == 1'd1) & (trunc_ln321_fu_726_p1 == 2'd2))) begin
            inputBuf_2_V_address1 = zext_ln202_fu_718_p1;
        end else if ((1'b1 == ap_condition_667)) begin
            inputBuf_2_V_address1 = zext_ln248_fu_606_p1;
        end else begin
            inputBuf_2_V_address1 = 'bx;
        end
    end else begin
        inputBuf_2_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_2_V_ce0 = 1'b1;
    end else begin
        inputBuf_2_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_2_V_ce1 = 1'b1;
    end else begin
        inputBuf_2_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_2_V_we1 = 1'b1;
    end else begin
        inputBuf_2_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_390_p2 == 1'd1) & (trunc_ln321_fu_726_p1 == 2'd3))) begin
            inputBuf_3_V_address1 = zext_ln202_fu_718_p1;
        end else if ((1'b1 == ap_condition_671)) begin
            inputBuf_3_V_address1 = zext_ln248_fu_606_p1;
        end else begin
            inputBuf_3_V_address1 = 'bx;
        end
    end else begin
        inputBuf_3_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_3_V_ce0 = 1'b1;
    end else begin
        inputBuf_3_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_3_V_ce1 = 1'b1;
    end else begin
        inputBuf_3_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_3_V_we1 = 1'b1;
    end else begin
        inputBuf_3_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln215_reg_891 == 1'd1) & (icmp_ln199_reg_887 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op205_write_state3 == 1'b1))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((icmp_ln197_fu_368_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((icmp_ln197_fu_368_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln197_fu_374_p2 = (i_0_0_reg_271 + 11'd1);

assign add_ln204_fu_730_p2 = (inp_15_0_fu_90 + 32'd1);

assign add_ln207_fu_746_p2 = (current_block_write_s_fu_106 + 32'd1);

assign add_ln211_fu_766_p2 = (read_block_1_0_fu_102 + 32'd1);

assign add_ln216_fu_421_p2 = (32'd1 + k_y_1_0_fu_86);

assign add_ln220_1_fu_453_p2 = (shl_ln_fu_445_p3 + count_simd_1_0_fu_98);

assign add_ln220_fu_439_p2 = (trunc_ln220_1_fu_435_p1 + trunc_ln220_fu_431_p1);

assign add_ln221_1_fu_467_p2 = (2'd1 + trunc_ln216_1_fu_427_p1);

assign add_ln221_fu_473_p2 = (add_ln221_1_fu_467_p2 + trunc_ln216_fu_417_p1);

assign add_ln223_fu_479_p2 = (32'd1 + count_simd_1_0_fu_98);

assign add_ln226_fu_496_p2 = (k_x_1_0_fu_94 + 32'd1);

assign add_ln232_fu_527_p2 = (ofm_x_1_0_fu_82 + 32'd1);

assign add_ln235_fu_547_p2 = (ofm_y_1_0_fu_78 + 32'd1);

assign add_ln256_1_fu_621_p2 = (trunc_ln197_fu_386_p1 + 2'd1);

assign add_ln256_fu_627_p2 = (current_block_write_s_fu_106 + 32'd1);

assign add_ln263_fu_693_p2 = (counter_internal_blo_fu_114 + 32'd1);

assign and_ln245_fu_600_p2 = (icmp_ln245_fu_588_p2 & icmp_ln245_1_fu_594_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

always @ (*) begin
    ap_block_pp0 = ((ap_ST_fsm_pp0_stage0 == ap_CS_fsm) & (1'b1 == ap_block_pp0_stage0_subdone));
end

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1)));
end

always @ (*) begin
    ap_block_state3_io = ((out_V_V_TREADY == 1'b0) & (ap_predicate_op205_write_state3 == 1'b1));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_230 = ((icmp_ln197_fu_368_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_condition_657 = ((1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd0));
end

always @ (*) begin
    ap_condition_663 = ((1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd1));
end

always @ (*) begin
    ap_condition_667 = ((1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd2));
end

always @ (*) begin
    ap_condition_671 = ((1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd3));
end

always @ (*) begin
    ap_enable_operation_127 = (ap_predicate_op127_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_129 = (ap_predicate_op129_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_131 = (ap_predicate_op131_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_133 = (ap_predicate_op133_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_170 = (ap_predicate_op170_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_172 = (ap_predicate_op172_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_174 = (ap_predicate_op174_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_176 = (ap_predicate_op176_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_200 = (ap_predicate_op200_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_201 = (ap_predicate_op201_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_202 = (ap_predicate_op202_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_203 = (ap_predicate_op203_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_65 = (ap_predicate_op65_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_67 = (ap_predicate_op67_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_69 = (ap_predicate_op69_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_71 = (ap_predicate_op71_load_state2 == 1'b1);
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

always @ (*) begin
    ap_enable_state2_pp0_iter0_stage0 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_enable_state3_pp0_iter1_stage0 = ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_predicate_op119_read_state2 = ((1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op127_store_state2 = ((1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd2));
end

always @ (*) begin
    ap_predicate_op129_store_state2 = ((1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd1));
end

always @ (*) begin
    ap_predicate_op131_store_state2 = ((1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd0));
end

always @ (*) begin
    ap_predicate_op133_store_state2 = ((1'd1 == and_ln245_fu_600_p2) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_1_fu_614_p1 == 2'd3));
end

always @ (*) begin
    ap_predicate_op162_read_state2 = ((icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op170_store_state2 = ((icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd2));
end

always @ (*) begin
    ap_predicate_op172_store_state2 = ((icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd1));
end

always @ (*) begin
    ap_predicate_op174_store_state2 = ((icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd0));
end

always @ (*) begin
    ap_predicate_op176_store_state2 = ((icmp_ln199_fu_390_p2 == 1'd1) & (icmp_ln197_fu_368_p2 == 1'd0) & (trunc_ln321_fu_726_p1 == 2'd3));
end

always @ (*) begin
    ap_predicate_op200_load_state3 = ((icmp_ln215_reg_891 == 1'd1) & (icmp_ln199_reg_887 == 1'd0));
end

always @ (*) begin
    ap_predicate_op201_load_state3 = ((icmp_ln215_reg_891 == 1'd1) & (icmp_ln199_reg_887 == 1'd0));
end

always @ (*) begin
    ap_predicate_op202_load_state3 = ((icmp_ln215_reg_891 == 1'd1) & (icmp_ln199_reg_887 == 1'd0));
end

always @ (*) begin
    ap_predicate_op203_load_state3 = ((icmp_ln215_reg_891 == 1'd1) & (icmp_ln199_reg_887 == 1'd0));
end

always @ (*) begin
    ap_predicate_op205_write_state3 = ((icmp_ln215_reg_891 == 1'd1) & (icmp_ln199_reg_887 == 1'd0));
end

always @ (*) begin
    ap_predicate_op65_load_state2 = ((icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op67_load_state2 = ((icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op69_load_state2 = ((icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op71_load_state2 = ((icmp_ln215_fu_399_p2 == 1'd1) & (icmp_ln199_fu_390_p2 == 1'd0) & (icmp_ln197_fu_368_p2 == 1'd0));
end

assign grp_fu_330_p2 = (current_line_1_0_fu_110 + 32'd1);

assign icmp_ln197_fu_368_p2 = ((i_0_0_reg_271 == 11'd1152) ? 1'b1 : 1'b0);

assign icmp_ln199_fu_390_p2 = ((inp_15_0_fu_90 < 32'd576) ? 1'b1 : 1'b0);

assign icmp_ln205_fu_342_p2 = ((grp_fu_330_p2 == 32'd192) ? 1'b1 : 1'b0);

assign icmp_ln208_fu_752_p2 = ((add_ln207_fu_746_p2 == 32'd4) ? 1'b1 : 1'b0);

assign icmp_ln215_fu_399_p2 = ((counter_internal_blo_fu_114 < 32'd575) ? 1'b1 : 1'b0);

assign icmp_ln224_fu_485_p2 = ((add_ln223_fu_479_p2 == 32'd64) ? 1'b1 : 1'b0);

assign icmp_ln227_fu_502_p2 = ((add_ln226_fu_496_p2 == 32'd3) ? 1'b1 : 1'b0);

assign icmp_ln230_fu_513_p2 = ((add_ln216_fu_421_p2 == 32'd3) ? 1'b1 : 1'b0);

assign icmp_ln233_fu_533_p2 = ((ofm_x_1_0_fu_82 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln236_fu_553_p2 = ((ofm_y_1_0_fu_78 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln245_1_fu_594_p2 = ((read_block_1_0_fu_102 < 32'd3) ? 1'b1 : 1'b0);

assign icmp_ln245_fu_588_p2 = ((counter_internal_blo_fu_114 < 32'd191) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_336_p2 = ((grp_fu_330_p2 == 32'd192) ? 1'b1 : 1'b0);

assign icmp_ln257_fu_633_p2 = ((add_ln256_fu_627_p2 == 32'd4) ? 1'b1 : 1'b0);

assign icmp_ln264_fu_699_p2 = ((add_ln263_fu_693_p2 == 32'd575) ? 1'b1 : 1'b0);

assign inputBuf_0_V_address0 = zext_ln221_fu_459_p1;

assign inputBuf_1_V_address0 = zext_ln221_fu_459_p1;

assign inputBuf_2_V_address0 = zext_ln221_fu_459_p1;

assign inputBuf_3_V_address0 = zext_ln221_fu_459_p1;

assign out_V_V_TDATA = tmp_V_1_fu_782_p6;

assign select_ln208_fu_758_p3 = ((icmp_ln208_fu_752_p2[0:0] === 1'b1) ? 32'd0 : add_ln207_fu_746_p2);

assign select_ln236_1_fu_567_p3 = ((icmp_ln236_fu_553_p2[0:0] === 1'b1) ? 32'd0 : add_ln235_fu_547_p2);

assign select_ln236_fu_559_p3 = ((icmp_ln236_fu_553_p2[0:0] === 1'b1) ? 32'd0 : inp_15_0_fu_90);

assign select_ln252_1_fu_655_p3 = ((icmp_ln252_fu_336_p2[0:0] === 1'b1) ? 32'd0 : grp_fu_330_p2);

assign select_ln252_2_fu_663_p3 = ((icmp_ln252_fu_336_p2[0:0] === 1'b1) ? add_ln256_1_fu_621_p2 : trunc_ln197_fu_386_p1);

assign select_ln252_fu_647_p3 = ((icmp_ln252_fu_336_p2[0:0] === 1'b1) ? select_ln257_fu_639_p3 : current_block_write_s_fu_106);

assign select_ln257_fu_639_p3 = ((icmp_ln257_fu_633_p2[0:0] === 1'b1) ? 32'd0 : add_ln256_fu_627_p2);

assign select_ln264_fu_705_p3 = ((icmp_ln264_fu_699_p2[0:0] === 1'b1) ? 32'd0 : add_ln263_fu_693_p2);

assign shl_ln_fu_445_p3 = {{add_ln220_fu_439_p2}, {6'd0}};

assign trunc_ln197_fu_386_p1 = read_block_1_0_fu_102[1:0];

assign trunc_ln216_1_fu_427_p1 = current_block_write_s_fu_106[1:0];

assign trunc_ln216_fu_417_p1 = k_y_1_0_fu_86[1:0];

assign trunc_ln220_1_fu_435_p1 = ofm_x_1_0_fu_82[25:0];

assign trunc_ln220_fu_431_p1 = k_x_1_0_fu_94[25:0];

assign trunc_ln321_1_fu_614_p1 = current_block_write_s_fu_106[1:0];

assign trunc_ln321_fu_726_p1 = current_block_write_s_fu_106[1:0];

assign zext_ln202_fu_718_p1 = current_line_1_0_fu_110;

assign zext_ln221_fu_459_p1 = add_ln220_1_fu_453_p2;

assign zext_ln248_fu_606_p1 = current_line_1_0_fu_110;

assign zext_ln252_fu_671_p1 = select_ln252_2_fu_663_p3;

endmodule //ConvolutionInputGenerator_1_ConvolutionInputGene_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbhl.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbhl_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbhl_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbhl(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbhl_rom Thresholding_Batch_0_Thresholding_Batcbhl_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actg8j.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actg8j_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actg8j_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actg8j(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actg8j_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actg8j_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actvdy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actvdy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actvdy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actvdy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actvdy_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actvdy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbfk.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbfk_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbfk_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbfk(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbfk_rom Thresholding_Batch_0_Thresholding_Batcbfk_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActqcK.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActqcK_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActqcK_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActqcK(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActqcK_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActqcK_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActwdI.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActwdI_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActwdI_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActwdI(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActwdI_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActwdI_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbgk.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbgk_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbgk_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbgk(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbgk_rom Thresholding_Batch_0_Thresholding_Batcbgk_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbkb_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 1;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbkb_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbkb(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd1;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbkb_rom Thresholding_Batch_0_Thresholding_Batcbkb_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batch_0.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="Thresholding_Batch_0_Thresholding_Batch_0,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=7.935000,HLS_SYN_LAT=3079,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=3467,HLS_SYN_LUT=6750,HLS_VERSION=2020_1_1}" *)

module Thresholding_Batch_0_Thresholding_Batch_0 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [7:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_Thresholding_Batch_fu_542_ap_start;
wire    grp_Thresholding_Batch_fu_542_ap_done;
wire    grp_Thresholding_Batch_fu_542_ap_idle;
wire    grp_Thresholding_Batch_fu_542_ap_ready;
wire    grp_Thresholding_Batch_fu_542_in_V_V_TREADY;
wire   [7:0] grp_Thresholding_Batch_fu_542_out_V_V_TDATA;
wire    grp_Thresholding_Batch_fu_542_out_V_V_TVALID;
wire    grp_Thresholding_Batch_fu_542_out_V_V_TREADY;
reg    grp_Thresholding_Batch_fu_542_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [7:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_Thresholding_Batch_fu_542_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

Thresholding_Batch_0_Thresholding_Batch grp_Thresholding_Batch_fu_542(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_Thresholding_Batch_fu_542_ap_start),
    .ap_done(grp_Thresholding_Batch_fu_542_ap_done),
    .ap_idle(grp_Thresholding_Batch_fu_542_ap_idle),
    .ap_ready(grp_Thresholding_Batch_fu_542_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_Thresholding_Batch_fu_542_in_V_V_TREADY),
    .out_V_V_TDATA(grp_Thresholding_Batch_fu_542_out_V_V_TDATA),
    .out_V_V_TVALID(grp_Thresholding_Batch_fu_542_out_V_V_TVALID),
    .out_V_V_TREADY(grp_Thresholding_Batch_fu_542_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_Thresholding_Batch_fu_542_out_V_V_TDATA),
    .vld_in(grp_Thresholding_Batch_fu_542_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_Thresholding_Batch_fu_542_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_Thresholding_Batch_fu_542_ap_start_reg <= 1'b1;
        end else if ((grp_Thresholding_Batch_fu_542_ap_ready == 1'b1)) begin
            grp_Thresholding_Batch_fu_542_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_Thresholding_Batch_fu_542_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_Thresholding_Batch_fu_542_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_Thresholding_Batch_fu_542_ap_start = grp_Thresholding_Batch_fu_542_ap_start_reg;

assign grp_Thresholding_Batch_fu_542_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //Thresholding_Batch_0_Thresholding_Batch_0
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_StreamingFCLayer_6jw.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

(* use_dsp = "no" *) module StreamingFCLayer_Batch_1_StreamingFCLayer_6jw_Mul_LUT_0(a, b, p);
input[4 - 1 : 0] a; 
input[4 - 1 : 0] b; 
output[8 - 1 : 0] p;

assign p = $signed(a) * $signed(b);
endmodule
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_StreamingFCLayer_6jw(
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



StreamingFCLayer_Batch_1_StreamingFCLayer_6jw_Mul_LUT_0 StreamingFCLayer_Batch_1_StreamingFCLayer_6jw_Mul_LUT_0_U(
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActOgC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActOgC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActOgC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActOgC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActOgC_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActOgC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/3a3d/hdl/verilog/StreamingDataWidthConverter_Batch_2_StreamingDataWidthCo_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingDataWidthConverter_Batch_2_StreamingDataWidthCo_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [15:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln402_fu_88_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln411_reg_154;
reg   [15:0] r_V_reg_61;
reg   [6:0] t_0_reg_72;
reg   [0:0] icmp_ln402_reg_135;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [6:0] t_fu_94_p2;
reg   [15:0] tmp_V_reg_144;
wire   [31:0] p_Result_s_fu_103_p3;
reg   [31:0] p_Result_s_reg_149;
wire   [0:0] icmp_ln411_fu_117_p2;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg   [15:0] ap_phi_mux_r_V_phi_fu_65_p4;
reg   [31:0] i_1_fu_44;
wire   [31:0] i_fu_111_p2;
reg    ap_block_pp0_stage0_01001;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_fu_117_p2 == 1'd0) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_1_fu_44 <= i_fu_111_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_fu_117_p2 == 1'd1) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        i_1_fu_44 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_reg_135 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        r_V_reg_61 <= tmp_V_reg_144;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        r_V_reg_61 <= 16'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        t_0_reg_72 <= t_fu_94_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        t_0_reg_72 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln402_reg_135 <= icmp_ln402_fu_88_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln411_reg_154 <= icmp_ln411_fu_117_p2;
        p_Result_s_reg_149 <= p_Result_s_fu_103_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_reg_144 <= in_V_V_TDATA;
    end
end

always @ (*) begin
    if ((icmp_ln402_fu_88_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln402_reg_135 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_r_V_phi_fu_65_p4 = tmp_V_reg_144;
    end else begin
        ap_phi_mux_r_V_phi_fu_65_p4 = r_V_reg_61;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln402_fu_88_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln411_reg_154 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_reg_154 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln402_fu_88_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln402_fu_88_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0));
end

always @ (*) begin
    ap_block_state3_io = ((icmp_ln411_reg_154 == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign i_fu_111_p2 = (i_1_fu_44 + 32'd1);

assign icmp_ln402_fu_88_p2 = ((t_0_reg_72 == 7'd64) ? 1'b1 : 1'b0);

assign icmp_ln411_fu_117_p2 = ((i_fu_111_p2 == 32'd2) ? 1'b1 : 1'b0);

assign out_V_V_TDATA = p_Result_s_reg_149;

assign p_Result_s_fu_103_p3 = {{in_V_V_TDATA}, {ap_phi_mux_r_V_phi_fu_65_p4}};

assign t_fu_94_p2 = (t_0_reg_72 + 7'd1);

endmodule //StreamingDataWidthConverter_Batch_2_StreamingDataWidthCo_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_8_0/synth/finn_design_StreamingFIFO_8_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_8:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_8,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_8_0,StreamingFIFO_8,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_8_0,StreamingFIFO_8,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_8,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_8_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [31 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 4, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [31 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 4, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_8 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActDeQ.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActDeQ_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActDeQ_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActDeQ(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActDeQ_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActDeQ_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ce70/StreamingFIFO_0.v


module StreamingFIFO_0(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [7:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(8)
)
StreamingFIFO_0_StreamingFIFO_0
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActRg6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActRg6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActRg6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActRg6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActRg6_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActRg6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcibs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_Batcibs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcibs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_Batcibs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_Batcibs_rom Thresholding_Batch_1_Thresholding_Batcibs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActpcA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActpcA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActpcA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActpcA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActpcA_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActpcA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActZio.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActZio_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActZio_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActZio(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActZio_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActZio_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_0_wstrm_0/synth/finn_design_StreamingFCLayer_Batch_0_wstrm_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:user:memstream:1.0
// IP Revision: 5

(* X_CORE_INFO = "memstream,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_0_wstrm_0,memstream,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_0_wstrm_0,memstream,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=user,x_ipName=memstream,x_ipVersion=1.0,x_ipCoreRevision=5,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED,CONFIG_EN=true,NSTREAMS=1,MEM_DEPTH=18432,MEM_WIDTH=32,MEM_INIT=/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_0_a2ilano3/,RAM_STYLE=auto,STRM0_WIDTH=32,STRM1_WIDTH=32,STRM2_WIDTH=32,STRM3_WIDTH=32,STRM4_WIDTH=32,STRM5_WIDTH=32,STR\
M0_DEPTH=18432,STRM1_DEPTH=2304,STRM2_DEPTH=2304,STRM3_DEPTH=2304,STRM4_DEPTH=2304,STRM5_DEPTH=2304,STRM0_OFFSET=0,STRM1_OFFSET=2304,STRM2_OFFSET=4608,STRM3_OFFSET=6912,STRM4_OFFSET=9216,STRM5_OFFSET=11520,AXILITE_ADDR_WIDTH=17}" *)
(* IP_DEFINITION_SOURCE = "package_project" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_0_wstrm_0 (
  aclk,
  aresetn,
  awready,
  awvalid,
  awaddr,
  awprot,
  wready,
  wvalid,
  wdata,
  wstrb,
  bready,
  bvalid,
  bresp,
  arready,
  arvalid,
  araddr,
  arprot,
  rready,
  rvalid,
  rresp,
  rdata,
  m_axis_0_tready,
  m_axis_0_tvalid,
  m_axis_0_tdata
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aclk, ASSOCIATED_BUSIF m_axis_0:m_axis_1:m_axis_2:m_axis_3:m_axis_4:m_axis_5:s_axilite, ASSOCIATED_RESET aresetn, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 aclk CLK" *)
input wire aclk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aresetn, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 aresetn RST" *)
input wire aresetn;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWREADY" *)
output wire awready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWVALID" *)
input wire awvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWADDR" *)
input wire [16 : 0] awaddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWPROT" *)
input wire [2 : 0] awprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WREADY" *)
output wire wready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WVALID" *)
input wire wvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WDATA" *)
input wire [31 : 0] wdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WSTRB" *)
input wire [3 : 0] wstrb;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BREADY" *)
input wire bready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BVALID" *)
output wire bvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BRESP" *)
output wire [1 : 0] bresp;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARREADY" *)
output wire arready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARVALID" *)
input wire arvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARADDR" *)
input wire [16 : 0] araddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARPROT" *)
input wire [2 : 0] arprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RREADY" *)
input wire rready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RVALID" *)
output wire rvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RRESP" *)
output wire [1 : 0] rresp;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axilite, DATA_WIDTH 32, PROTOCOL AXI4LITE, FREQ_HZ 100000000.000000, ID_WIDTH 0, ADDR_WIDTH 17, AWUSER_WIDTH 0, ARUSER_WIDTH 0, WUSER_WIDTH 0, RUSER_WIDTH 0, BUSER_WIDTH 0, READ_WRITE_MODE READ_WRITE, HAS_BURST 0, HAS_LOCK 0, HAS_PROT 1, HAS_CACHE 0, HAS_QOS 0, HAS_REGION 0, HAS_WSTRB 1, HAS_BRESP 1, HAS_RRESP 1, SUPPORTS_NARROW_BURST 0, NUM_READ_OUTSTANDING 1, NUM_WRITE_OUTSTANDING 1, MAX_BURST_LENGTH 1, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, NUM_READ_THREADS 1, NUM_W\
RITE_THREADS 1, RUSER_BITS_PER_BYTE 0, WUSER_BITS_PER_BYTE 0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RDATA" *)
output wire [31 : 0] rdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TREADY" *)
input wire m_axis_0_tready;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TVALID" *)
output wire m_axis_0_tvalid;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME m_axis_0, TDATA_NUM_BYTES 4, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TDATA" *)
output wire [31 : 0] m_axis_0_tdata;

  memstream #(
    .CONFIG_EN(1'B1),
    .NSTREAMS(1),
    .MEM_DEPTH(18432),
    .MEM_WIDTH(32),
    .MEM_INIT("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_0_a2ilano3/"),
    .RAM_STYLE("auto"),
    .STRM0_WIDTH(32),
    .STRM1_WIDTH(32),
    .STRM2_WIDTH(32),
    .STRM3_WIDTH(32),
    .STRM4_WIDTH(32),
    .STRM5_WIDTH(32),
    .STRM0_DEPTH(18432),
    .STRM1_DEPTH(2304),
    .STRM2_DEPTH(2304),
    .STRM3_DEPTH(2304),
    .STRM4_DEPTH(2304),
    .STRM5_DEPTH(2304),
    .STRM0_OFFSET(0),
    .STRM1_OFFSET(2304),
    .STRM2_OFFSET(4608),
    .STRM3_OFFSET(6912),
    .STRM4_OFFSET(9216),
    .STRM5_OFFSET(11520),
    .AXILITE_ADDR_WIDTH(17)
  ) inst (
    .aclk(aclk),
    .aresetn(aresetn),
    .awready(awready),
    .awvalid(awvalid),
    .awaddr(awaddr),
    .awprot(awprot),
    .wready(wready),
    .wvalid(wvalid),
    .wdata(wdata),
    .wstrb(wstrb),
    .bready(bready),
    .bvalid(bvalid),
    .bresp(bresp),
    .arready(arready),
    .arvalid(arvalid),
    .araddr(araddr),
    .arprot(arprot),
    .rready(rready),
    .rvalid(rvalid),
    .rresp(rresp),
    .rdata(rdata),
    .m_axis_0_afull(1'B0),
    .m_axis_0_tready(m_axis_0_tready),
    .m_axis_0_tvalid(m_axis_0_tvalid),
    .m_axis_0_tdata(m_axis_0_tdata),
    .m_axis_1_afull(1'B0),
    .m_axis_1_tready(1'B1),
    .m_axis_1_tvalid(),
    .m_axis_1_tdata(),
    .m_axis_2_afull(1'B0),
    .m_axis_2_tready(1'B1),
    .m_axis_2_tvalid(),
    .m_axis_2_tdata(),
    .m_axis_3_afull(1'B0),
    .m_axis_3_tready(1'B1),
    .m_axis_3_tvalid(),
    .m_axis_3_tdata(),
    .m_axis_4_afull(1'B0),
    .m_axis_4_tready(1'B1),
    .m_axis_4_tvalid(),
    .m_axis_4_tdata(),
    .m_axis_5_afull(1'B0),
    .m_axis_5_tready(1'B1),
    .m_axis_5_tvalid(),
    .m_axis_5_tdata()
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbzo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbzo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbzo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbzo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbzo_rom Thresholding_Batch_0_Thresholding_Batcbzo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actudo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actudo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actudo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actudo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actudo_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actudo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccNA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccNA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccNA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccNA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccNA_rom Thresholding_Batch_0_Thresholding_BatccNA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActAem.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActAem_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActAem_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActAem(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActAem_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActAem_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actibs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actibs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actibs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actibs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actibs_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actibs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActThq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActThq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActThq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActThq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActThq_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActThq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActeOg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActeOg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActeOg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActeOg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActeOg_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActeOg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActIfE.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActIfE_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActIfE_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActIfE(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActIfE_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActIfE_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/abe7/hdl/verilog/ConvolutionInputGenerator_0_ConvolutionInputGene_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module ConvolutionInputGenerator_0_ConvolutionInputGene_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [7:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln197_fu_374_p2;
wire   [0:0] icmp_ln199_fu_396_p2;
wire   [0:0] and_ln245_fu_606_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln199_reg_893;
reg   [0:0] icmp_ln215_reg_897;
reg   [15:0] i_0_0_reg_277;
reg    ap_predicate_op119_read_state2;
reg    ap_predicate_op162_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_predicate_op205_write_state3;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [15:0] add_ln197_fu_380_p2;
wire   [0:0] icmp_ln215_fu_405_p2;
wire   [1:0] add_ln221_fu_479_p2;
reg   [1:0] add_ln221_reg_901;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
wire   [9:0] inputBuf_0_V_address0;
reg    inputBuf_0_V_ce0;
wire   [7:0] inputBuf_0_V_q0;
reg   [9:0] inputBuf_0_V_address1;
reg    inputBuf_0_V_ce1;
reg    inputBuf_0_V_we1;
wire   [9:0] inputBuf_1_V_address0;
reg    inputBuf_1_V_ce0;
wire   [7:0] inputBuf_1_V_q0;
reg   [9:0] inputBuf_1_V_address1;
reg    inputBuf_1_V_ce1;
reg    inputBuf_1_V_we1;
wire   [9:0] inputBuf_2_V_address0;
reg    inputBuf_2_V_ce0;
wire   [7:0] inputBuf_2_V_q0;
reg   [9:0] inputBuf_2_V_address1;
reg    inputBuf_2_V_ce1;
reg    inputBuf_2_V_we1;
wire   [9:0] inputBuf_3_V_address0;
reg    inputBuf_3_V_ce0;
wire   [7:0] inputBuf_3_V_q0;
reg   [9:0] inputBuf_3_V_address1;
reg    inputBuf_3_V_ce1;
reg    inputBuf_3_V_we1;
wire   [63:0] zext_ln221_fu_465_p1;
wire   [63:0] zext_ln248_fu_612_p1;
wire   [63:0] zext_ln202_fu_724_p1;
reg   [31:0] ofm_y_1_0_fu_84;
wire   [31:0] select_ln236_1_fu_573_p3;
wire   [0:0] icmp_ln224_fu_491_p2;
wire   [0:0] icmp_ln227_fu_508_p2;
wire   [0:0] icmp_ln230_fu_519_p2;
wire   [0:0] icmp_ln233_fu_539_p2;
reg   [31:0] ofm_x_1_0_fu_88;
wire   [31:0] add_ln232_fu_533_p2;
reg   [31:0] k_y_1_0_fu_92;
wire   [31:0] add_ln216_fu_427_p2;
reg   [31:0] inp_15_0_fu_96;
wire   [31:0] select_ln236_fu_565_p3;
wire   [31:0] add_ln204_fu_736_p2;
reg   [31:0] k_x_1_0_fu_100;
wire   [31:0] add_ln226_fu_502_p2;
reg   [31:0] count_simd_1_0_fu_104;
wire   [31:0] add_ln223_fu_485_p2;
reg   [31:0] read_block_1_0_fu_108;
wire   [31:0] zext_ln252_fu_677_p1;
wire   [31:0] add_ln211_fu_772_p2;
wire   [0:0] icmp_ln205_fu_348_p2;
reg   [31:0] current_block_write_s_fu_112;
wire   [31:0] select_ln252_fu_653_p3;
wire   [31:0] select_ln208_fu_764_p3;
reg   [31:0] current_line_1_0_fu_116;
wire   [31:0] select_ln252_1_fu_661_p3;
wire   [31:0] grp_fu_336_p2;
reg   [31:0] counter_internal_blo_fu_120;
wire   [31:0] select_ln264_fu_711_p3;
wire   [7:0] tmp_V_1_fu_788_p6;
reg    ap_block_pp0_stage0_01001;
wire   [1:0] trunc_ln321_1_fu_620_p1;
wire   [1:0] trunc_ln321_fu_732_p1;
wire   [25:0] trunc_ln220_1_fu_441_p1;
wire   [25:0] trunc_ln220_fu_437_p1;
wire   [25:0] add_ln220_fu_445_p2;
wire   [31:0] shl_ln_fu_451_p3;
wire   [31:0] add_ln220_1_fu_459_p2;
wire   [1:0] trunc_ln216_1_fu_433_p1;
wire   [1:0] add_ln221_1_fu_473_p2;
wire   [1:0] trunc_ln216_fu_423_p1;
wire   [31:0] add_ln235_fu_553_p2;
wire   [0:0] icmp_ln236_fu_559_p2;
wire   [0:0] icmp_ln245_fu_594_p2;
wire   [0:0] icmp_ln245_1_fu_600_p2;
wire   [3:0] trunc_ln197_fu_392_p1;
wire   [31:0] add_ln256_fu_633_p2;
wire   [0:0] icmp_ln257_fu_639_p2;
wire   [0:0] icmp_ln252_fu_342_p2;
wire   [31:0] select_ln257_fu_645_p3;
wire   [3:0] add_ln256_1_fu_627_p2;
wire   [3:0] select_ln252_2_fu_669_p3;
wire   [31:0] add_ln263_fu_699_p2;
wire   [0:0] icmp_ln264_fu_705_p2;
wire   [31:0] add_ln207_fu_752_p2;
wire   [0:0] icmp_ln208_fu_758_p2;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_block_pp0;
reg    ap_predicate_op127_store_state2;
reg    ap_enable_operation_127;
reg    ap_enable_state2_pp0_iter0_stage0;
reg    ap_predicate_op69_load_state2;
reg    ap_enable_operation_69;
reg    ap_predicate_op202_load_state3;
reg    ap_enable_operation_202;
reg    ap_enable_state3_pp0_iter1_stage0;
reg    ap_predicate_op170_store_state2;
reg    ap_enable_operation_170;
reg    ap_predicate_op129_store_state2;
reg    ap_enable_operation_129;
reg    ap_predicate_op67_load_state2;
reg    ap_enable_operation_67;
reg    ap_predicate_op201_load_state3;
reg    ap_enable_operation_201;
reg    ap_predicate_op172_store_state2;
reg    ap_enable_operation_172;
reg    ap_predicate_op131_store_state2;
reg    ap_enable_operation_131;
reg    ap_predicate_op65_load_state2;
reg    ap_enable_operation_65;
reg    ap_predicate_op200_load_state3;
reg    ap_enable_operation_200;
reg    ap_predicate_op174_store_state2;
reg    ap_enable_operation_174;
reg    ap_predicate_op133_store_state2;
reg    ap_enable_operation_133;
reg    ap_predicate_op71_load_state2;
reg    ap_enable_operation_71;
reg    ap_predicate_op203_load_state3;
reg    ap_enable_operation_203;
reg    ap_predicate_op176_store_state2;
reg    ap_enable_operation_176;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_660;
reg    ap_condition_230;
reg    ap_condition_666;
reg    ap_condition_670;
reg    ap_condition_674;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

ConvolutionInputGenerator_0_ConvolutionInputGbkb #(
    .DataWidth( 8 ),
    .AddressRange( 768 ),
    .AddressWidth( 10 ))
inputBuf_0_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_0_V_address0),
    .ce0(inputBuf_0_V_ce0),
    .q0(inputBuf_0_V_q0),
    .address1(inputBuf_0_V_address1),
    .ce1(inputBuf_0_V_ce1),
    .we1(inputBuf_0_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_0_ConvolutionInputGbkb #(
    .DataWidth( 8 ),
    .AddressRange( 768 ),
    .AddressWidth( 10 ))
inputBuf_1_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_1_V_address0),
    .ce0(inputBuf_1_V_ce0),
    .q0(inputBuf_1_V_q0),
    .address1(inputBuf_1_V_address1),
    .ce1(inputBuf_1_V_ce1),
    .we1(inputBuf_1_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_0_ConvolutionInputGbkb #(
    .DataWidth( 8 ),
    .AddressRange( 768 ),
    .AddressWidth( 10 ))
inputBuf_2_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_2_V_address0),
    .ce0(inputBuf_2_V_ce0),
    .q0(inputBuf_2_V_q0),
    .address1(inputBuf_2_V_address1),
    .ce1(inputBuf_2_V_ce1),
    .we1(inputBuf_2_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_0_ConvolutionInputGbkb #(
    .DataWidth( 8 ),
    .AddressRange( 768 ),
    .AddressWidth( 10 ))
inputBuf_3_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(inputBuf_3_V_address0),
    .ce0(inputBuf_3_V_ce0),
    .q0(inputBuf_3_V_q0),
    .address1(inputBuf_3_V_address1),
    .ce1(inputBuf_3_V_ce1),
    .we1(inputBuf_3_V_we1),
    .d1(in_V_V_TDATA)
);

ConvolutionInputGenerator_0_ConvolutionInputGfYi #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 8 ),
    .din1_WIDTH( 8 ),
    .din2_WIDTH( 8 ),
    .din3_WIDTH( 8 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 8 ))
ConvolutionInputGfYi_U1(
    .din0(inputBuf_0_V_q0),
    .din1(inputBuf_1_V_q0),
    .din2(inputBuf_2_V_q0),
    .din3(inputBuf_3_V_q0),
    .din4(add_ln221_reg_901),
    .dout(tmp_V_1_fu_788_p6)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln224_fu_491_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        count_simd_1_0_fu_104 <= add_ln223_fu_485_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln227_fu_508_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln230_fu_519_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln233_fu_539_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln233_fu_539_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        count_simd_1_0_fu_104 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        counter_internal_blo_fu_120 <= select_ln264_fu_711_p3;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_348_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        counter_internal_blo_fu_120 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_348_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_block_write_s_fu_112 <= select_ln208_fu_764_p3;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_block_write_s_fu_112 <= select_ln252_fu_653_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        current_block_write_s_fu_112 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln205_fu_348_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_line_1_0_fu_116 <= grp_fu_336_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        current_line_1_0_fu_116 <= select_ln252_1_fu_661_p3;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_348_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        current_line_1_0_fu_116 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_0_reg_277 <= 16'd0;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_0_reg_277 <= add_ln197_fu_380_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inp_15_0_fu_96 <= add_ln204_fu_736_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln233_fu_539_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inp_15_0_fu_96 <= select_ln236_fu_565_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        inp_15_0_fu_96 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln227_fu_508_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        k_x_1_0_fu_100 <= add_ln226_fu_502_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln230_fu_519_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln233_fu_539_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln233_fu_539_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        k_x_1_0_fu_100 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln230_fu_519_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        k_y_1_0_fu_92 <= add_ln216_fu_427_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        k_y_1_0_fu_92 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln233_fu_539_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ofm_x_1_0_fu_88 <= add_ln232_fu_533_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln233_fu_539_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ofm_x_1_0_fu_88 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln233_fu_539_p2 == 1'd1) & (icmp_ln230_fu_519_p2 == 1'd1) & (icmp_ln227_fu_508_p2 == 1'd1) & (icmp_ln224_fu_491_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ofm_y_1_0_fu_84 <= select_ln236_1_fu_573_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        ofm_y_1_0_fu_84 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln205_fu_348_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        read_block_1_0_fu_108 <= add_ln211_fu_772_p2;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        read_block_1_0_fu_108 <= zext_ln252_fu_677_p1;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        read_block_1_0_fu_108 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln221_reg_901 <= add_ln221_fu_479_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln197_fu_374_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln199_reg_893 <= icmp_ln199_fu_396_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln215_reg_897 <= icmp_ln215_fu_405_p2;
    end
end

always @ (*) begin
    if ((icmp_ln197_fu_374_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op119_read_state2 == 1'b1)))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_396_p2 == 1'd1) & (trunc_ln321_fu_732_p1 == 2'd0))) begin
            inputBuf_0_V_address1 = zext_ln202_fu_724_p1;
        end else if ((1'b1 == ap_condition_660)) begin
            inputBuf_0_V_address1 = zext_ln248_fu_612_p1;
        end else begin
            inputBuf_0_V_address1 = 'bx;
        end
    end else begin
        inputBuf_0_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_0_V_ce0 = 1'b1;
    end else begin
        inputBuf_0_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_0_V_ce1 = 1'b1;
    end else begin
        inputBuf_0_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_0_V_we1 = 1'b1;
    end else begin
        inputBuf_0_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_396_p2 == 1'd1) & (trunc_ln321_fu_732_p1 == 2'd1))) begin
            inputBuf_1_V_address1 = zext_ln202_fu_724_p1;
        end else if ((1'b1 == ap_condition_666)) begin
            inputBuf_1_V_address1 = zext_ln248_fu_612_p1;
        end else begin
            inputBuf_1_V_address1 = 'bx;
        end
    end else begin
        inputBuf_1_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_1_V_ce0 = 1'b1;
    end else begin
        inputBuf_1_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_1_V_ce1 = 1'b1;
    end else begin
        inputBuf_1_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_1_V_we1 = 1'b1;
    end else begin
        inputBuf_1_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_396_p2 == 1'd1) & (trunc_ln321_fu_732_p1 == 2'd2))) begin
            inputBuf_2_V_address1 = zext_ln202_fu_724_p1;
        end else if ((1'b1 == ap_condition_670)) begin
            inputBuf_2_V_address1 = zext_ln248_fu_612_p1;
        end else begin
            inputBuf_2_V_address1 = 'bx;
        end
    end else begin
        inputBuf_2_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_2_V_ce0 = 1'b1;
    end else begin
        inputBuf_2_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_2_V_ce1 = 1'b1;
    end else begin
        inputBuf_2_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_2_V_we1 = 1'b1;
    end else begin
        inputBuf_2_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_condition_230)) begin
        if (((icmp_ln199_fu_396_p2 == 1'd1) & (trunc_ln321_fu_732_p1 == 2'd3))) begin
            inputBuf_3_V_address1 = zext_ln202_fu_724_p1;
        end else if ((1'b1 == ap_condition_674)) begin
            inputBuf_3_V_address1 = zext_ln248_fu_612_p1;
        end else begin
            inputBuf_3_V_address1 = 'bx;
        end
    end else begin
        inputBuf_3_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        inputBuf_3_V_ce0 = 1'b1;
    end else begin
        inputBuf_3_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_3_V_ce1 = 1'b1;
    end else begin
        inputBuf_3_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        inputBuf_3_V_we1 = 1'b1;
    end else begin
        inputBuf_3_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op205_write_state3 == 1'b1))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((icmp_ln197_fu_374_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((icmp_ln197_fu_374_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln197_fu_380_p2 = (i_0_0_reg_277 + 16'd1);

assign add_ln204_fu_736_p2 = (inp_15_0_fu_96 + 32'd1);

assign add_ln207_fu_752_p2 = (current_block_write_s_fu_112 + 32'd1);

assign add_ln211_fu_772_p2 = (read_block_1_0_fu_108 + 32'd1);

assign add_ln216_fu_427_p2 = (32'd1 + k_y_1_0_fu_92);

assign add_ln220_1_fu_459_p2 = (shl_ln_fu_451_p3 + count_simd_1_0_fu_104);

assign add_ln220_fu_445_p2 = (trunc_ln220_1_fu_441_p1 + trunc_ln220_fu_437_p1);

assign add_ln221_1_fu_473_p2 = (2'd1 + trunc_ln216_1_fu_433_p1);

assign add_ln221_fu_479_p2 = (add_ln221_1_fu_473_p2 + trunc_ln216_fu_423_p1);

assign add_ln223_fu_485_p2 = (32'd1 + count_simd_1_0_fu_104);

assign add_ln226_fu_502_p2 = (k_x_1_0_fu_100 + 32'd1);

assign add_ln232_fu_533_p2 = (ofm_x_1_0_fu_88 + 32'd1);

assign add_ln235_fu_553_p2 = (ofm_y_1_0_fu_84 + 32'd1);

assign add_ln256_1_fu_627_p2 = (trunc_ln197_fu_392_p1 + 4'd1);

assign add_ln256_fu_633_p2 = (current_block_write_s_fu_112 + 32'd1);

assign add_ln263_fu_699_p2 = (counter_internal_blo_fu_120 + 32'd1);

assign and_ln245_fu_606_p2 = (icmp_ln245_fu_594_p2 & icmp_ln245_1_fu_600_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

always @ (*) begin
    ap_block_pp0 = ((ap_ST_fsm_pp0_stage0 == ap_CS_fsm) & (1'b1 == ap_block_pp0_stage0_subdone));
end

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((in_V_V_TVALID == 1'b0) & (ap_predicate_op119_read_state2 == 1'b1)));
end

always @ (*) begin
    ap_block_state3_io = ((out_V_V_TREADY == 1'b0) & (ap_predicate_op205_write_state3 == 1'b1));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_230 = ((icmp_ln197_fu_374_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_condition_660 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd0));
end

always @ (*) begin
    ap_condition_666 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd1));
end

always @ (*) begin
    ap_condition_670 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd2));
end

always @ (*) begin
    ap_condition_674 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd3));
end

always @ (*) begin
    ap_enable_operation_127 = (ap_predicate_op127_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_129 = (ap_predicate_op129_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_131 = (ap_predicate_op131_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_133 = (ap_predicate_op133_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_170 = (ap_predicate_op170_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_172 = (ap_predicate_op172_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_174 = (ap_predicate_op174_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_176 = (ap_predicate_op176_store_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_200 = (ap_predicate_op200_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_201 = (ap_predicate_op201_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_202 = (ap_predicate_op202_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_203 = (ap_predicate_op203_load_state3 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_65 = (ap_predicate_op65_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_67 = (ap_predicate_op67_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_69 = (ap_predicate_op69_load_state2 == 1'b1);
end

always @ (*) begin
    ap_enable_operation_71 = (ap_predicate_op71_load_state2 == 1'b1);
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

always @ (*) begin
    ap_enable_state2_pp0_iter0_stage0 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_enable_state3_pp0_iter1_stage0 = ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

always @ (*) begin
    ap_predicate_op119_read_state2 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op127_store_state2 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd2));
end

always @ (*) begin
    ap_predicate_op129_store_state2 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd1));
end

always @ (*) begin
    ap_predicate_op131_store_state2 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd0));
end

always @ (*) begin
    ap_predicate_op133_store_state2 = ((1'd1 == and_ln245_fu_606_p2) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_1_fu_620_p1 == 2'd3));
end

always @ (*) begin
    ap_predicate_op162_read_state2 = ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op170_store_state2 = ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd2));
end

always @ (*) begin
    ap_predicate_op172_store_state2 = ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd1));
end

always @ (*) begin
    ap_predicate_op174_store_state2 = ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd0));
end

always @ (*) begin
    ap_predicate_op176_store_state2 = ((icmp_ln199_fu_396_p2 == 1'd1) & (icmp_ln197_fu_374_p2 == 1'd0) & (trunc_ln321_fu_732_p1 == 2'd3));
end

always @ (*) begin
    ap_predicate_op200_load_state3 = ((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0));
end

always @ (*) begin
    ap_predicate_op201_load_state3 = ((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0));
end

always @ (*) begin
    ap_predicate_op202_load_state3 = ((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0));
end

always @ (*) begin
    ap_predicate_op203_load_state3 = ((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0));
end

always @ (*) begin
    ap_predicate_op205_write_state3 = ((icmp_ln215_reg_897 == 1'd1) & (icmp_ln199_reg_893 == 1'd0));
end

always @ (*) begin
    ap_predicate_op65_load_state2 = ((icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op67_load_state2 = ((icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op69_load_state2 = ((icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0));
end

always @ (*) begin
    ap_predicate_op71_load_state2 = ((icmp_ln215_fu_405_p2 == 1'd1) & (icmp_ln199_fu_396_p2 == 1'd0) & (icmp_ln197_fu_374_p2 == 1'd0));
end

assign grp_fu_336_p2 = (current_line_1_0_fu_116 + 32'd1);

assign icmp_ln197_fu_374_p2 = ((i_0_0_reg_277 == 16'd59904) ? 1'b1 : 1'b0);

assign icmp_ln199_fu_396_p2 = ((inp_15_0_fu_96 < 32'd2304) ? 1'b1 : 1'b0);

assign icmp_ln205_fu_348_p2 = ((grp_fu_336_p2 == 32'd768) ? 1'b1 : 1'b0);

assign icmp_ln208_fu_758_p2 = ((add_ln207_fu_752_p2 == 32'd4) ? 1'b1 : 1'b0);

assign icmp_ln215_fu_405_p2 = ((counter_internal_blo_fu_120 < 32'd5759) ? 1'b1 : 1'b0);

assign icmp_ln224_fu_491_p2 = ((add_ln223_fu_485_p2 == 32'd64) ? 1'b1 : 1'b0);

assign icmp_ln227_fu_508_p2 = ((add_ln226_fu_502_p2 == 32'd3) ? 1'b1 : 1'b0);

assign icmp_ln230_fu_519_p2 = ((add_ln216_fu_427_p2 == 32'd3) ? 1'b1 : 1'b0);

assign icmp_ln233_fu_539_p2 = ((add_ln232_fu_533_p2 == 32'd10) ? 1'b1 : 1'b0);

assign icmp_ln236_fu_559_p2 = ((add_ln235_fu_553_p2 == 32'd10) ? 1'b1 : 1'b0);

assign icmp_ln245_1_fu_600_p2 = ((read_block_1_0_fu_108 < 32'd12) ? 1'b1 : 1'b0);

assign icmp_ln245_fu_594_p2 = ((counter_internal_blo_fu_120 < 32'd767) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_342_p2 = ((grp_fu_336_p2 == 32'd768) ? 1'b1 : 1'b0);

assign icmp_ln257_fu_639_p2 = ((add_ln256_fu_633_p2 == 32'd4) ? 1'b1 : 1'b0);

assign icmp_ln264_fu_705_p2 = ((add_ln263_fu_699_p2 == 32'd5759) ? 1'b1 : 1'b0);

assign inputBuf_0_V_address0 = zext_ln221_fu_465_p1;

assign inputBuf_1_V_address0 = zext_ln221_fu_465_p1;

assign inputBuf_2_V_address0 = zext_ln221_fu_465_p1;

assign inputBuf_3_V_address0 = zext_ln221_fu_465_p1;

assign out_V_V_TDATA = tmp_V_1_fu_788_p6;

assign select_ln208_fu_764_p3 = ((icmp_ln208_fu_758_p2[0:0] === 1'b1) ? 32'd0 : add_ln207_fu_752_p2);

assign select_ln236_1_fu_573_p3 = ((icmp_ln236_fu_559_p2[0:0] === 1'b1) ? 32'd0 : add_ln235_fu_553_p2);

assign select_ln236_fu_565_p3 = ((icmp_ln236_fu_559_p2[0:0] === 1'b1) ? 32'd0 : inp_15_0_fu_96);

assign select_ln252_1_fu_661_p3 = ((icmp_ln252_fu_342_p2[0:0] === 1'b1) ? 32'd0 : grp_fu_336_p2);

assign select_ln252_2_fu_669_p3 = ((icmp_ln252_fu_342_p2[0:0] === 1'b1) ? add_ln256_1_fu_627_p2 : trunc_ln197_fu_392_p1);

assign select_ln252_fu_653_p3 = ((icmp_ln252_fu_342_p2[0:0] === 1'b1) ? select_ln257_fu_645_p3 : current_block_write_s_fu_112);

assign select_ln257_fu_645_p3 = ((icmp_ln257_fu_639_p2[0:0] === 1'b1) ? 32'd0 : add_ln256_fu_633_p2);

assign select_ln264_fu_711_p3 = ((icmp_ln264_fu_705_p2[0:0] === 1'b1) ? 32'd0 : add_ln263_fu_699_p2);

assign shl_ln_fu_451_p3 = {{add_ln220_fu_445_p2}, {6'd0}};

assign trunc_ln197_fu_392_p1 = read_block_1_0_fu_108[3:0];

assign trunc_ln216_1_fu_433_p1 = current_block_write_s_fu_112[1:0];

assign trunc_ln216_fu_423_p1 = k_y_1_0_fu_92[1:0];

assign trunc_ln220_1_fu_441_p1 = ofm_x_1_0_fu_88[25:0];

assign trunc_ln220_fu_437_p1 = k_x_1_0_fu_100[25:0];

assign trunc_ln321_1_fu_620_p1 = current_block_write_s_fu_112[1:0];

assign trunc_ln321_fu_732_p1 = current_block_write_s_fu_112[1:0];

assign zext_ln202_fu_724_p1 = current_line_1_0_fu_116;

assign zext_ln221_fu_465_p1 = add_ln220_1_fu_459_p2;

assign zext_ln248_fu_612_p1 = current_line_1_0_fu_116;

assign zext_ln252_fu_677_p1 = select_ln252_2_fu_669_p3;

endmodule //ConvolutionInputGenerator_0_ConvolutionInputGene_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actbkb_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actbkb_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actbkb(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actbkb_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actbkb_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccPA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccPA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccPA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccPA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccPA_rom Thresholding_Batch_0_Thresholding_BatccPA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbkl.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbkl_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbkl_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbkl(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbkl_rom Thresholding_Batch_0_Thresholding_Batcbkl_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_5_wstrm_0/synth/finn_design_StreamingFCLayer_Batch_5_wstrm_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:user:memstream:1.0
// IP Revision: 5

(* X_CORE_INFO = "memstream,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_5_wstrm_0,memstream,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_5_wstrm_0,memstream,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=user,x_ipName=memstream,x_ipVersion=1.0,x_ipCoreRevision=5,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED,CONFIG_EN=true,NSTREAMS=1,MEM_DEPTH=4608,MEM_WIDTH=32,MEM_INIT=/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_5_g5ap2jtp/,RAM_STYLE=auto,STRM0_WIDTH=32,STRM1_WIDTH=32,STRM2_WIDTH=32,STRM3_WIDTH=32,STRM4_WIDTH=32,STRM5_WIDTH=32,STRM\
0_DEPTH=4608,STRM1_DEPTH=2304,STRM2_DEPTH=2304,STRM3_DEPTH=2304,STRM4_DEPTH=2304,STRM5_DEPTH=2304,STRM0_OFFSET=0,STRM1_OFFSET=2304,STRM2_OFFSET=4608,STRM3_OFFSET=6912,STRM4_OFFSET=9216,STRM5_OFFSET=11520,AXILITE_ADDR_WIDTH=15}" *)
(* IP_DEFINITION_SOURCE = "package_project" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_5_wstrm_0 (
  aclk,
  aresetn,
  awready,
  awvalid,
  awaddr,
  awprot,
  wready,
  wvalid,
  wdata,
  wstrb,
  bready,
  bvalid,
  bresp,
  arready,
  arvalid,
  araddr,
  arprot,
  rready,
  rvalid,
  rresp,
  rdata,
  m_axis_0_tready,
  m_axis_0_tvalid,
  m_axis_0_tdata
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aclk, ASSOCIATED_BUSIF m_axis_0:m_axis_1:m_axis_2:m_axis_3:m_axis_4:m_axis_5:s_axilite, ASSOCIATED_RESET aresetn, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 aclk CLK" *)
input wire aclk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aresetn, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 aresetn RST" *)
input wire aresetn;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWREADY" *)
output wire awready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWVALID" *)
input wire awvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWADDR" *)
input wire [14 : 0] awaddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWPROT" *)
input wire [2 : 0] awprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WREADY" *)
output wire wready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WVALID" *)
input wire wvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WDATA" *)
input wire [31 : 0] wdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WSTRB" *)
input wire [3 : 0] wstrb;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BREADY" *)
input wire bready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BVALID" *)
output wire bvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BRESP" *)
output wire [1 : 0] bresp;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARREADY" *)
output wire arready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARVALID" *)
input wire arvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARADDR" *)
input wire [14 : 0] araddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARPROT" *)
input wire [2 : 0] arprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RREADY" *)
input wire rready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RVALID" *)
output wire rvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RRESP" *)
output wire [1 : 0] rresp;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axilite, DATA_WIDTH 32, PROTOCOL AXI4LITE, FREQ_HZ 100000000.000000, ID_WIDTH 0, ADDR_WIDTH 15, AWUSER_WIDTH 0, ARUSER_WIDTH 0, WUSER_WIDTH 0, RUSER_WIDTH 0, BUSER_WIDTH 0, READ_WRITE_MODE READ_WRITE, HAS_BURST 0, HAS_LOCK 0, HAS_PROT 1, HAS_CACHE 0, HAS_QOS 0, HAS_REGION 0, HAS_WSTRB 1, HAS_BRESP 1, HAS_RRESP 1, SUPPORTS_NARROW_BURST 0, NUM_READ_OUTSTANDING 1, NUM_WRITE_OUTSTANDING 1, MAX_BURST_LENGTH 1, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, NUM_READ_THREADS 1, NUM_W\
RITE_THREADS 1, RUSER_BITS_PER_BYTE 0, WUSER_BITS_PER_BYTE 0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RDATA" *)
output wire [31 : 0] rdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TREADY" *)
input wire m_axis_0_tready;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TVALID" *)
output wire m_axis_0_tvalid;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME m_axis_0, TDATA_NUM_BYTES 4, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TDATA" *)
output wire [31 : 0] m_axis_0_tdata;

  memstream #(
    .CONFIG_EN(1'B1),
    .NSTREAMS(1),
    .MEM_DEPTH(4608),
    .MEM_WIDTH(32),
    .MEM_INIT("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_5_g5ap2jtp/"),
    .RAM_STYLE("auto"),
    .STRM0_WIDTH(32),
    .STRM1_WIDTH(32),
    .STRM2_WIDTH(32),
    .STRM3_WIDTH(32),
    .STRM4_WIDTH(32),
    .STRM5_WIDTH(32),
    .STRM0_DEPTH(4608),
    .STRM1_DEPTH(2304),
    .STRM2_DEPTH(2304),
    .STRM3_DEPTH(2304),
    .STRM4_DEPTH(2304),
    .STRM5_DEPTH(2304),
    .STRM0_OFFSET(0),
    .STRM1_OFFSET(2304),
    .STRM2_OFFSET(4608),
    .STRM3_OFFSET(6912),
    .STRM4_OFFSET(9216),
    .STRM5_OFFSET(11520),
    .AXILITE_ADDR_WIDTH(15)
  ) inst (
    .aclk(aclk),
    .aresetn(aresetn),
    .awready(awready),
    .awvalid(awvalid),
    .awaddr(awaddr),
    .awprot(awprot),
    .wready(wready),
    .wvalid(wvalid),
    .wdata(wdata),
    .wstrb(wstrb),
    .bready(bready),
    .bvalid(bvalid),
    .bresp(bresp),
    .arready(arready),
    .arvalid(arvalid),
    .araddr(araddr),
    .arprot(arprot),
    .rready(rready),
    .rvalid(rvalid),
    .rresp(rresp),
    .rdata(rdata),
    .m_axis_0_afull(1'B0),
    .m_axis_0_tready(m_axis_0_tready),
    .m_axis_0_tvalid(m_axis_0_tvalid),
    .m_axis_0_tdata(m_axis_0_tdata),
    .m_axis_1_afull(1'B0),
    .m_axis_1_tready(1'B1),
    .m_axis_1_tvalid(),
    .m_axis_1_tdata(),
    .m_axis_2_afull(1'B0),
    .m_axis_2_tready(1'B1),
    .m_axis_2_tvalid(),
    .m_axis_2_tdata(),
    .m_axis_3_afull(1'B0),
    .m_axis_3_tready(1'B1),
    .m_axis_3_tvalid(),
    .m_axis_3_tdata(),
    .m_axis_4_afull(1'B0),
    .m_axis_4_tready(1'B1),
    .m_axis_4_tvalid(),
    .m_axis_4_tdata(),
    .m_axis_5_afull(1'B0),
    .m_axis_5_tready(1'B1),
    .m_axis_5_tvalid(),
    .m_axis_5_tdata()
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/5192/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcibs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_Batcibs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcibs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_Batcibs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_Batcibs_rom Thresholding_Batch_2_Thresholding_Batcibs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Activa.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingFCLayer_Batch_3_Matrix_Vector_Activa (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY,
        weight_V_V_TDATA,
        weight_V_V_TVALID,
        weight_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state7 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [31:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;
input  [127:0] weight_V_V_TDATA;
input   weight_V_V_TVALID;
output   weight_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;
reg weight_V_V_TREADY;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [6:0] threshs_m_thresholds_55_address0;
reg    threshs_m_thresholds_55_ce0;
wire   [14:0] threshs_m_thresholds_55_q0;
wire   [6:0] threshs_m_thresholds_54_address0;
reg    threshs_m_thresholds_54_ce0;
wire   [14:0] threshs_m_thresholds_54_q0;
wire   [6:0] threshs_m_thresholds_49_address0;
reg    threshs_m_thresholds_49_ce0;
wire   [15:0] threshs_m_thresholds_49_q0;
wire   [6:0] threshs_m_thresholds_48_address0;
reg    threshs_m_thresholds_48_ce0;
wire   [15:0] threshs_m_thresholds_48_q0;
wire   [6:0] threshs_m_thresholds_47_address0;
reg    threshs_m_thresholds_47_ce0;
wire   [15:0] threshs_m_thresholds_47_q0;
wire   [6:0] threshs_m_thresholds_46_address0;
reg    threshs_m_thresholds_46_ce0;
wire   [15:0] threshs_m_thresholds_46_q0;
wire   [6:0] threshs_m_thresholds_45_address0;
reg    threshs_m_thresholds_45_ce0;
wire   [15:0] threshs_m_thresholds_45_q0;
wire   [6:0] threshs_m_thresholds_44_address0;
reg    threshs_m_thresholds_44_ce0;
wire   [15:0] threshs_m_thresholds_44_q0;
wire   [6:0] threshs_m_thresholds_43_address0;
reg    threshs_m_thresholds_43_ce0;
wire   [15:0] threshs_m_thresholds_43_q0;
wire   [6:0] threshs_m_thresholds_42_address0;
reg    threshs_m_thresholds_42_ce0;
wire   [15:0] threshs_m_thresholds_42_q0;
wire   [6:0] threshs_m_thresholds_53_address0;
reg    threshs_m_thresholds_53_ce0;
wire   [15:0] threshs_m_thresholds_53_q0;
wire   [6:0] threshs_m_thresholds_52_address0;
reg    threshs_m_thresholds_52_ce0;
wire   [15:0] threshs_m_thresholds_52_q0;
wire   [6:0] threshs_m_thresholds_51_address0;
reg    threshs_m_thresholds_51_ce0;
wire   [15:0] threshs_m_thresholds_51_q0;
wire   [6:0] threshs_m_thresholds_50_address0;
reg    threshs_m_thresholds_50_ce0;
wire   [15:0] threshs_m_thresholds_50_q0;
wire   [6:0] threshs_m_thresholds_41_address0;
reg    threshs_m_thresholds_41_ce0;
wire   [15:0] threshs_m_thresholds_41_q0;
wire   [6:0] threshs_m_thresholds_40_address0;
reg    threshs_m_thresholds_40_ce0;
wire   [15:0] threshs_m_thresholds_40_q0;
wire   [6:0] threshs_m_thresholds_35_address0;
reg    threshs_m_thresholds_35_ce0;
wire   [15:0] threshs_m_thresholds_35_q0;
wire   [6:0] threshs_m_thresholds_34_address0;
reg    threshs_m_thresholds_34_ce0;
wire   [15:0] threshs_m_thresholds_34_q0;
wire   [6:0] threshs_m_thresholds_33_address0;
reg    threshs_m_thresholds_33_ce0;
wire   [14:0] threshs_m_thresholds_33_q0;
wire   [6:0] threshs_m_thresholds_32_address0;
reg    threshs_m_thresholds_32_ce0;
wire   [14:0] threshs_m_thresholds_32_q0;
wire   [6:0] threshs_m_thresholds_31_address0;
reg    threshs_m_thresholds_31_ce0;
wire   [14:0] threshs_m_thresholds_31_q0;
wire   [6:0] threshs_m_thresholds_30_address0;
reg    threshs_m_thresholds_30_ce0;
wire   [14:0] threshs_m_thresholds_30_q0;
wire   [6:0] threshs_m_thresholds_29_address0;
reg    threshs_m_thresholds_29_ce0;
wire   [14:0] threshs_m_thresholds_29_q0;
wire   [6:0] threshs_m_thresholds_28_address0;
reg    threshs_m_thresholds_28_ce0;
wire   [14:0] threshs_m_thresholds_28_q0;
wire   [6:0] threshs_m_thresholds_39_address0;
reg    threshs_m_thresholds_39_ce0;
wire   [14:0] threshs_m_thresholds_39_q0;
wire   [6:0] threshs_m_thresholds_38_address0;
reg    threshs_m_thresholds_38_ce0;
wire   [14:0] threshs_m_thresholds_38_q0;
wire   [6:0] threshs_m_thresholds_37_address0;
reg    threshs_m_thresholds_37_ce0;
wire   [14:0] threshs_m_thresholds_37_q0;
wire   [6:0] threshs_m_thresholds_36_address0;
reg    threshs_m_thresholds_36_ce0;
wire   [14:0] threshs_m_thresholds_36_q0;
wire   [6:0] threshs_m_thresholds_27_address0;
reg    threshs_m_thresholds_27_ce0;
wire   [15:0] threshs_m_thresholds_27_q0;
wire   [6:0] threshs_m_thresholds_26_address0;
reg    threshs_m_thresholds_26_ce0;
wire   [15:0] threshs_m_thresholds_26_q0;
wire   [6:0] threshs_m_thresholds_21_address0;
reg    threshs_m_thresholds_21_ce0;
wire   [15:0] threshs_m_thresholds_21_q0;
wire   [6:0] threshs_m_thresholds_20_address0;
reg    threshs_m_thresholds_20_ce0;
wire   [15:0] threshs_m_thresholds_20_q0;
wire   [6:0] threshs_m_thresholds_19_address0;
reg    threshs_m_thresholds_19_ce0;
wire   [15:0] threshs_m_thresholds_19_q0;
wire   [6:0] threshs_m_thresholds_18_address0;
reg    threshs_m_thresholds_18_ce0;
wire   [15:0] threshs_m_thresholds_18_q0;
wire   [6:0] threshs_m_thresholds_17_address0;
reg    threshs_m_thresholds_17_ce0;
wire   [15:0] threshs_m_thresholds_17_q0;
wire   [6:0] threshs_m_thresholds_16_address0;
reg    threshs_m_thresholds_16_ce0;
wire   [15:0] threshs_m_thresholds_16_q0;
wire   [6:0] threshs_m_thresholds_15_address0;
reg    threshs_m_thresholds_15_ce0;
wire   [15:0] threshs_m_thresholds_15_q0;
wire   [6:0] threshs_m_thresholds_14_address0;
reg    threshs_m_thresholds_14_ce0;
wire   [15:0] threshs_m_thresholds_14_q0;
wire   [6:0] threshs_m_thresholds_25_address0;
reg    threshs_m_thresholds_25_ce0;
wire   [15:0] threshs_m_thresholds_25_q0;
wire   [6:0] threshs_m_thresholds_24_address0;
reg    threshs_m_thresholds_24_ce0;
wire   [15:0] threshs_m_thresholds_24_q0;
wire   [6:0] threshs_m_thresholds_23_address0;
reg    threshs_m_thresholds_23_ce0;
wire   [15:0] threshs_m_thresholds_23_q0;
wire   [6:0] threshs_m_thresholds_22_address0;
reg    threshs_m_thresholds_22_ce0;
wire   [15:0] threshs_m_thresholds_22_q0;
wire   [6:0] threshs_m_thresholds_13_address0;
reg    threshs_m_thresholds_13_ce0;
wire   [15:0] threshs_m_thresholds_13_q0;
wire   [6:0] threshs_m_thresholds_12_address0;
reg    threshs_m_thresholds_12_ce0;
wire   [15:0] threshs_m_thresholds_12_q0;
wire   [6:0] threshs_m_thresholds_7_address0;
reg    threshs_m_thresholds_7_ce0;
wire   [15:0] threshs_m_thresholds_7_q0;
wire   [6:0] threshs_m_thresholds_6_address0;
reg    threshs_m_thresholds_6_ce0;
wire   [15:0] threshs_m_thresholds_6_q0;
wire   [6:0] threshs_m_thresholds_5_address0;
reg    threshs_m_thresholds_5_ce0;
wire   [15:0] threshs_m_thresholds_5_q0;
wire   [6:0] threshs_m_thresholds_4_address0;
reg    threshs_m_thresholds_4_ce0;
wire   [15:0] threshs_m_thresholds_4_q0;
wire   [6:0] threshs_m_thresholds_3_address0;
reg    threshs_m_thresholds_3_ce0;
wire   [15:0] threshs_m_thresholds_3_q0;
wire   [6:0] threshs_m_thresholds_2_address0;
reg    threshs_m_thresholds_2_ce0;
wire   [15:0] threshs_m_thresholds_2_q0;
wire   [6:0] threshs_m_thresholds_1_address0;
reg    threshs_m_thresholds_1_ce0;
wire   [15:0] threshs_m_thresholds_1_q0;
wire   [6:0] threshs_m_thresholds_address0;
reg    threshs_m_thresholds_ce0;
wire   [15:0] threshs_m_thresholds_q0;
wire   [6:0] threshs_m_thresholds_11_address0;
reg    threshs_m_thresholds_11_ce0;
wire   [15:0] threshs_m_thresholds_11_q0;
wire   [6:0] threshs_m_thresholds_10_address0;
reg    threshs_m_thresholds_10_ce0;
wire   [15:0] threshs_m_thresholds_10_q0;
wire   [6:0] threshs_m_thresholds_9_address0;
reg    threshs_m_thresholds_9_ce0;
wire   [15:0] threshs_m_thresholds_9_q0;
wire   [6:0] threshs_m_thresholds_8_address0;
reg    threshs_m_thresholds_8_ce0;
wire   [15:0] threshs_m_thresholds_8_q0;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln248_fu_1359_p2;
wire   [0:0] icmp_ln252_fu_1374_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter4;
reg   [0:0] icmp_ln289_reg_4790;
reg   [0:0] icmp_ln289_reg_4790_pp0_iter3_reg;
reg    weight_V_V_TDATA_blk_n;
reg   [12:0] i_0_reg_1267;
reg    ap_predicate_op98_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
reg    ap_block_state6_io;
reg    ap_block_pp0_stage0_11001;
wire   [12:0] i_fu_1365_p2;
wire   [31:0] inElem_V_1_fu_1483_p34;
wire   [4:0] trunc_ln321_fu_1553_p1;
wire   [0:0] icmp_ln271_fu_1720_p2;
reg   [0:0] icmp_ln271_reg_4622;
reg   [0:0] icmp_ln271_reg_4622_pp0_iter1_reg;
wire   [3:0] wgt_M_instance_0_V_fu_1726_p1;
reg  signed [3:0] wgt_M_instance_0_V_reg_4630;
reg  signed [3:0] wgt_M_instance_1_V_reg_4635;
reg  signed [3:0] wgt_M_instance_2_V_reg_4640;
reg  signed [3:0] wgt_M_instance_3_V_reg_4645;
reg  signed [3:0] wgt_M_instance_4_V_reg_4650;
reg  signed [3:0] wgt_M_instance_5_V_reg_4655;
reg  signed [3:0] wgt_M_instance_6_V_reg_4660;
reg  signed [3:0] wgt_M_instance_7_V_reg_4665;
reg  signed [3:0] wgt_M_instance_0_V_1_reg_4670;
reg  signed [3:0] wgt_M_instance_1_V_1_reg_4675;
reg  signed [3:0] wgt_M_instance_2_V_1_reg_4680;
reg  signed [3:0] wgt_M_instance_3_V_1_reg_4685;
reg  signed [3:0] wgt_M_instance_4_V_1_reg_4690;
reg  signed [3:0] wgt_M_instance_5_V_1_reg_4695;
reg  signed [3:0] wgt_M_instance_6_V_1_reg_4700;
reg  signed [3:0] wgt_M_instance_7_V_1_reg_4705;
reg  signed [3:0] wgt_M_instance_0_V_2_reg_4710;
reg  signed [3:0] wgt_M_instance_1_V_2_reg_4715;
reg  signed [3:0] wgt_M_instance_2_V_2_reg_4720;
reg  signed [3:0] wgt_M_instance_3_V_2_reg_4725;
reg  signed [3:0] wgt_M_instance_4_V_2_reg_4730;
reg  signed [3:0] wgt_M_instance_5_V_2_reg_4735;
reg  signed [3:0] wgt_M_instance_6_V_2_reg_4740;
reg  signed [3:0] wgt_M_instance_7_V_2_reg_4745;
reg  signed [3:0] wgt_M_instance_0_V_3_reg_4750;
reg  signed [3:0] wgt_M_instance_1_V_3_reg_4755;
reg  signed [3:0] wgt_M_instance_2_V_3_reg_4760;
reg  signed [3:0] wgt_M_instance_3_V_3_reg_4765;
reg  signed [3:0] wgt_M_instance_4_V_3_reg_4770;
reg  signed [3:0] wgt_M_instance_5_V_3_reg_4775;
reg  signed [3:0] wgt_M_instance_6_V_3_reg_4780;
reg  signed [3:0] wgt_M_instance_7_V_3_reg_4785;
wire   [0:0] icmp_ln289_fu_2046_p2;
reg   [0:0] icmp_ln289_reg_4790_pp0_iter1_reg;
reg   [0:0] icmp_ln289_reg_4790_pp0_iter2_reg;
wire  signed [7:0] mul_ln1352_5_fu_2203_p2;
reg  signed [7:0] mul_ln1352_5_reg_4794;
wire   [8:0] add_ln700_1_fu_2263_p2;
reg   [8:0] add_ln700_1_reg_4799;
wire   [8:0] add_ln700_3_fu_2269_p2;
reg   [8:0] add_ln700_3_reg_4804;
wire   [9:0] add_ln700_5_fu_2285_p2;
reg   [9:0] add_ln700_5_reg_4809;
wire  signed [7:0] mul_ln1352_13_fu_2359_p2;
reg  signed [7:0] mul_ln1352_13_reg_4814;
wire   [8:0] add_ln700_9_fu_2391_p2;
reg   [8:0] add_ln700_9_reg_4819;
wire   [8:0] add_ln700_11_fu_2397_p2;
reg   [8:0] add_ln700_11_reg_4824;
wire   [9:0] add_ln700_13_fu_2413_p2;
reg   [9:0] add_ln700_13_reg_4829;
wire  signed [7:0] mul_ln1352_21_fu_2487_p2;
reg  signed [7:0] mul_ln1352_21_reg_4834;
wire   [8:0] add_ln700_17_fu_2519_p2;
reg   [8:0] add_ln700_17_reg_4839;
wire   [8:0] add_ln700_19_fu_2525_p2;
reg   [8:0] add_ln700_19_reg_4844;
wire   [9:0] add_ln700_21_fu_2541_p2;
reg   [9:0] add_ln700_21_reg_4849;
wire  signed [7:0] mul_ln1352_29_fu_2615_p2;
reg  signed [7:0] mul_ln1352_29_reg_4854;
wire   [8:0] add_ln700_25_fu_2647_p2;
reg   [8:0] add_ln700_25_reg_4859;
wire   [8:0] add_ln700_27_fu_2653_p2;
reg   [8:0] add_ln700_27_reg_4864;
wire   [9:0] add_ln700_29_fu_2669_p2;
reg   [9:0] add_ln700_29_reg_4869;
wire   [0:0] icmp_ln899_fu_2987_p2;
reg   [0:0] icmp_ln899_reg_5154;
reg   [0:0] icmp_ln899_reg_5154_pp0_iter3_reg;
wire   [0:0] icmp_ln899_1_fu_2997_p2;
reg   [0:0] icmp_ln899_1_reg_5159;
reg   [0:0] icmp_ln899_1_reg_5159_pp0_iter3_reg;
wire   [0:0] icmp_ln899_2_fu_3003_p2;
reg   [0:0] icmp_ln899_2_reg_5164;
reg   [0:0] icmp_ln899_2_reg_5164_pp0_iter3_reg;
wire   [0:0] icmp_ln899_3_fu_3009_p2;
reg   [0:0] icmp_ln899_3_reg_5169;
wire   [0:0] icmp_ln899_4_fu_3015_p2;
reg   [0:0] icmp_ln899_4_reg_5174;
wire   [0:0] icmp_ln899_5_fu_3021_p2;
reg   [0:0] icmp_ln899_5_reg_5179;
wire   [0:0] icmp_ln899_6_fu_3027_p2;
reg   [0:0] icmp_ln899_6_reg_5184;
wire   [0:0] icmp_ln899_7_fu_3033_p2;
reg   [0:0] icmp_ln899_7_reg_5189;
wire   [0:0] icmp_ln899_8_fu_3039_p2;
reg   [0:0] icmp_ln899_8_reg_5194;
wire   [0:0] icmp_ln899_9_fu_3045_p2;
reg   [0:0] icmp_ln899_9_reg_5199;
wire   [0:0] icmp_ln899_10_fu_3051_p2;
reg   [0:0] icmp_ln899_10_reg_5204;
wire   [0:0] icmp_ln899_11_fu_3057_p2;
reg   [0:0] icmp_ln899_11_reg_5209;
wire   [0:0] icmp_ln899_12_fu_3063_p2;
reg   [0:0] icmp_ln899_12_reg_5214;
wire   [0:0] icmp_ln899_13_fu_3069_p2;
reg   [0:0] icmp_ln899_13_reg_5219;
wire   [0:0] icmp_ln899_14_fu_3075_p2;
reg   [0:0] icmp_ln899_14_reg_5224;
reg   [0:0] icmp_ln899_14_reg_5224_pp0_iter3_reg;
wire   [0:0] icmp_ln899_15_fu_3081_p2;
reg   [0:0] icmp_ln899_15_reg_5229;
reg   [0:0] icmp_ln899_15_reg_5229_pp0_iter3_reg;
wire   [0:0] icmp_ln899_16_fu_3087_p2;
reg   [0:0] icmp_ln899_16_reg_5234;
reg   [0:0] icmp_ln899_16_reg_5234_pp0_iter3_reg;
wire   [0:0] icmp_ln899_17_fu_3093_p2;
reg   [0:0] icmp_ln899_17_reg_5239;
wire   [0:0] icmp_ln899_18_fu_3103_p2;
reg   [0:0] icmp_ln899_18_reg_5244;
wire   [0:0] icmp_ln899_19_fu_3113_p2;
reg   [0:0] icmp_ln899_19_reg_5249;
wire   [0:0] icmp_ln899_20_fu_3123_p2;
reg   [0:0] icmp_ln899_20_reg_5254;
wire   [0:0] icmp_ln899_21_fu_3133_p2;
reg   [0:0] icmp_ln899_21_reg_5259;
wire   [0:0] icmp_ln899_22_fu_3143_p2;
reg   [0:0] icmp_ln899_22_reg_5264;
wire   [0:0] icmp_ln899_23_fu_3153_p2;
reg   [0:0] icmp_ln899_23_reg_5269;
wire   [0:0] icmp_ln899_24_fu_3163_p2;
reg   [0:0] icmp_ln899_24_reg_5274;
wire   [0:0] icmp_ln899_25_fu_3173_p2;
reg   [0:0] icmp_ln899_25_reg_5279;
wire   [0:0] icmp_ln899_26_fu_3183_p2;
reg   [0:0] icmp_ln899_26_reg_5284;
wire   [0:0] icmp_ln899_27_fu_3193_p2;
reg   [0:0] icmp_ln899_27_reg_5289;
wire   [0:0] icmp_ln899_28_fu_3199_p2;
reg   [0:0] icmp_ln899_28_reg_5294;
reg   [0:0] icmp_ln899_28_reg_5294_pp0_iter3_reg;
wire   [0:0] icmp_ln899_29_fu_3205_p2;
reg   [0:0] icmp_ln899_29_reg_5299;
reg   [0:0] icmp_ln899_29_reg_5299_pp0_iter3_reg;
wire   [0:0] icmp_ln899_30_fu_3211_p2;
reg   [0:0] icmp_ln899_30_reg_5304;
reg   [0:0] icmp_ln899_30_reg_5304_pp0_iter3_reg;
wire   [0:0] icmp_ln899_31_fu_3217_p2;
reg   [0:0] icmp_ln899_31_reg_5309;
wire   [0:0] icmp_ln899_32_fu_3223_p2;
reg   [0:0] icmp_ln899_32_reg_5314;
wire   [0:0] icmp_ln899_33_fu_3229_p2;
reg   [0:0] icmp_ln899_33_reg_5319;
wire   [0:0] icmp_ln899_34_fu_3235_p2;
reg   [0:0] icmp_ln899_34_reg_5324;
wire   [0:0] icmp_ln899_35_fu_3241_p2;
reg   [0:0] icmp_ln899_35_reg_5329;
wire   [0:0] icmp_ln899_36_fu_3247_p2;
reg   [0:0] icmp_ln899_36_reg_5334;
wire   [0:0] icmp_ln899_37_fu_3253_p2;
reg   [0:0] icmp_ln899_37_reg_5339;
wire   [0:0] icmp_ln899_38_fu_3259_p2;
reg   [0:0] icmp_ln899_38_reg_5344;
wire   [0:0] icmp_ln899_39_fu_3265_p2;
reg   [0:0] icmp_ln899_39_reg_5349;
wire   [0:0] icmp_ln899_40_fu_3271_p2;
reg   [0:0] icmp_ln899_40_reg_5354;
wire   [0:0] icmp_ln899_41_fu_3277_p2;
reg   [0:0] icmp_ln899_41_reg_5359;
wire   [0:0] icmp_ln899_42_fu_3283_p2;
reg   [0:0] icmp_ln899_42_reg_5364;
reg   [0:0] icmp_ln899_42_reg_5364_pp0_iter3_reg;
wire   [0:0] icmp_ln899_43_fu_3289_p2;
reg   [0:0] icmp_ln899_43_reg_5369;
reg   [0:0] icmp_ln899_43_reg_5369_pp0_iter3_reg;
wire   [0:0] icmp_ln899_44_fu_3295_p2;
reg   [0:0] icmp_ln899_44_reg_5374;
reg   [0:0] icmp_ln899_44_reg_5374_pp0_iter3_reg;
wire   [0:0] icmp_ln899_45_fu_3301_p2;
reg   [0:0] icmp_ln899_45_reg_5379;
wire   [0:0] icmp_ln899_46_fu_3307_p2;
reg   [0:0] icmp_ln899_46_reg_5384;
wire   [0:0] icmp_ln899_47_fu_3313_p2;
reg   [0:0] icmp_ln899_47_reg_5389;
wire   [0:0] icmp_ln899_48_fu_3319_p2;
reg   [0:0] icmp_ln899_48_reg_5394;
wire   [0:0] icmp_ln899_49_fu_3325_p2;
reg   [0:0] icmp_ln899_49_reg_5399;
wire   [0:0] icmp_ln899_50_fu_3331_p2;
reg   [0:0] icmp_ln899_50_reg_5404;
wire   [0:0] icmp_ln899_51_fu_3337_p2;
reg   [0:0] icmp_ln899_51_reg_5409;
wire   [0:0] icmp_ln899_52_fu_3343_p2;
reg   [0:0] icmp_ln899_52_reg_5414;
wire   [0:0] icmp_ln899_53_fu_3349_p2;
reg   [0:0] icmp_ln899_53_reg_5419;
wire   [0:0] icmp_ln899_54_fu_3355_p2;
reg   [0:0] icmp_ln899_54_reg_5424;
wire   [0:0] icmp_ln899_55_fu_3361_p2;
reg   [0:0] icmp_ln899_55_reg_5429;
wire   [2:0] add_ln700_36_fu_3486_p2;
reg   [2:0] add_ln700_36_reg_5434;
wire   [2:0] add_ln700_43_fu_3534_p2;
reg   [2:0] add_ln700_43_reg_5439;
wire   [2:0] add_ln700_49_fu_3659_p2;
reg   [2:0] add_ln700_49_reg_5444;
wire   [2:0] add_ln700_56_fu_3707_p2;
reg   [2:0] add_ln700_56_reg_5449;
wire   [2:0] add_ln700_62_fu_3832_p2;
reg   [2:0] add_ln700_62_reg_5454;
wire   [2:0] add_ln700_69_fu_3880_p2;
reg   [2:0] add_ln700_69_reg_5459;
wire   [2:0] add_ln700_75_fu_4005_p2;
reg   [2:0] add_ln700_75_reg_5464;
wire   [2:0] add_ln700_82_fu_4053_p2;
reg   [2:0] add_ln700_82_reg_5469;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
wire   [31:0] ap_phi_reg_pp0_iter0_act_m_val_V_reg_1278;
reg   [31:0] ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278;
wire   [63:0] zext_ln142_fu_2678_p1;
reg   [15:0] accu_V_0_0_0_fu_368;
wire   [15:0] accu_0_0_V_fu_2837_p2;
reg   [15:0] accu_V_0_1_0_fu_372;
wire   [15:0] accu_0_1_V_fu_2877_p2;
reg   [15:0] accu_V_0_2_0_fu_376;
wire   [15:0] accu_0_2_V_fu_2917_p2;
reg   [15:0] accu_V_0_3_0_fu_380;
wire   [15:0] accu_0_3_V_fu_2957_p2;
reg   [31:0] sf_1_fu_384;
wire   [31:0] sf_fu_2040_p2;
reg   [31:0] tmp_V_fu_388;
reg   [31:0] tmp_V_1_fu_392;
reg   [31:0] tmp_V_2_fu_396;
reg   [31:0] tmp_V_4_fu_400;
reg   [31:0] tmp_V_5_fu_404;
reg   [31:0] tmp_V_6_fu_408;
reg   [31:0] tmp_V_7_fu_412;
reg   [31:0] tmp_V_8_fu_416;
reg   [31:0] tmp_V_9_fu_420;
reg   [31:0] tmp_V_10_fu_424;
reg   [31:0] tmp_V_11_fu_428;
reg   [31:0] tmp_V_12_fu_432;
reg   [31:0] tmp_V_13_fu_436;
reg   [31:0] tmp_V_14_fu_440;
reg   [31:0] tmp_V_15_fu_444;
reg   [31:0] tmp_V_16_fu_448;
reg   [31:0] tmp_V_17_fu_452;
reg   [31:0] tmp_V_18_fu_456;
reg   [31:0] tmp_V_19_fu_460;
reg   [31:0] tmp_V_20_fu_464;
reg   [31:0] tmp_V_21_fu_468;
reg   [31:0] tmp_V_22_fu_472;
reg   [31:0] tmp_V_23_fu_476;
reg   [31:0] tmp_V_24_fu_480;
reg   [31:0] tmp_V_25_fu_484;
reg   [31:0] tmp_V_26_fu_488;
reg   [31:0] tmp_V_27_fu_492;
reg   [31:0] tmp_V_28_fu_496;
reg   [31:0] tmp_V_29_fu_500;
reg   [31:0] tmp_V_30_fu_504;
reg   [31:0] tmp_V_31_fu_508;
reg   [31:0] tmp_V_32_fu_512;
reg   [31:0] nf_assign_fu_516;
wire   [31:0] select_ln301_fu_2750_p3;
reg   [31:0] ap_sig_allocacmp_nf_assign_load_1;
reg    ap_block_pp0_stage0_01001;
wire   [4:0] inElem_V_1_fu_1483_p33;
wire   [3:0] trunc_ln647_fu_2057_p1;
wire   [3:0] mul_ln1352_fu_2068_p0;
wire   [7:0] zext_ln215_fu_2064_p1;
wire  signed [7:0] mul_ln1352_fu_2068_p2;
wire   [3:0] arg_V_read_assign_1_fu_2078_p4;
wire   [3:0] mul_ln1352_1_fu_2095_p0;
wire   [7:0] zext_ln215_1_fu_2091_p1;
wire  signed [7:0] mul_ln1352_1_fu_2095_p2;
wire   [3:0] arg_V_read_assign_2_fu_2105_p4;
wire   [3:0] mul_ln1352_2_fu_2122_p0;
wire   [7:0] zext_ln215_2_fu_2118_p1;
wire  signed [7:0] mul_ln1352_2_fu_2122_p2;
wire   [3:0] arg_V_read_assign_3_fu_2132_p4;
wire   [3:0] mul_ln1352_3_fu_2149_p0;
wire   [7:0] zext_ln215_3_fu_2145_p1;
wire  signed [7:0] mul_ln1352_3_fu_2149_p2;
wire   [3:0] arg_V_read_assign_4_fu_2159_p4;
wire   [3:0] mul_ln1352_4_fu_2176_p0;
wire   [7:0] zext_ln215_4_fu_2172_p1;
wire  signed [7:0] mul_ln1352_4_fu_2176_p2;
wire   [3:0] arg_V_read_assign_5_fu_2186_p4;
wire   [3:0] mul_ln1352_5_fu_2203_p0;
wire   [7:0] zext_ln215_5_fu_2199_p1;
wire   [3:0] arg_V_read_assign_6_fu_2209_p4;
wire   [3:0] mul_ln1352_6_fu_2226_p0;
wire   [7:0] zext_ln215_6_fu_2222_p1;
wire  signed [7:0] mul_ln1352_6_fu_2226_p2;
wire   [3:0] arg_V_read_assign_7_fu_2236_p4;
wire   [3:0] mul_ln1352_7_fu_2253_p0;
wire   [7:0] zext_ln215_7_fu_2249_p1;
wire  signed [7:0] mul_ln1352_7_fu_2253_p2;
wire  signed [8:0] sext_ln170_4_fu_2182_p1;
wire  signed [8:0] sext_ln170_5_fu_2232_p1;
wire  signed [8:0] sext_ln170_fu_2074_p1;
wire  signed [8:0] sext_ln170_3_fu_2155_p1;
wire  signed [8:0] sext_ln700_1_fu_2259_p1;
wire  signed [8:0] sext_ln170_1_fu_2101_p1;
wire   [8:0] add_ln700_4_fu_2275_p2;
wire  signed [9:0] sext_ln170_2_fu_2128_p1;
wire  signed [9:0] sext_ln700_4_fu_2281_p1;
wire   [3:0] mul_ln1352_8_fu_2294_p0;
wire  signed [7:0] mul_ln1352_8_fu_2294_p2;
wire   [3:0] mul_ln1352_9_fu_2307_p0;
wire  signed [7:0] mul_ln1352_9_fu_2307_p2;
wire   [3:0] mul_ln1352_10_fu_2320_p0;
wire  signed [7:0] mul_ln1352_10_fu_2320_p2;
wire   [3:0] mul_ln1352_11_fu_2333_p0;
wire  signed [7:0] mul_ln1352_11_fu_2333_p2;
wire   [3:0] mul_ln1352_12_fu_2346_p0;
wire  signed [7:0] mul_ln1352_12_fu_2346_p2;
wire   [3:0] mul_ln1352_13_fu_2359_p0;
wire   [3:0] mul_ln1352_14_fu_2368_p0;
wire  signed [7:0] mul_ln1352_14_fu_2368_p2;
wire   [3:0] mul_ln1352_15_fu_2381_p0;
wire  signed [7:0] mul_ln1352_15_fu_2381_p2;
wire  signed [8:0] sext_ln170_10_fu_2352_p1;
wire  signed [8:0] sext_ln170_11_fu_2374_p1;
wire  signed [8:0] sext_ln170_6_fu_2300_p1;
wire  signed [8:0] sext_ln170_9_fu_2339_p1;
wire  signed [8:0] sext_ln700_8_fu_2387_p1;
wire  signed [8:0] sext_ln170_7_fu_2313_p1;
wire   [8:0] add_ln700_12_fu_2403_p2;
wire  signed [9:0] sext_ln170_8_fu_2326_p1;
wire  signed [9:0] sext_ln700_11_fu_2409_p1;
wire   [3:0] mul_ln1352_16_fu_2422_p0;
wire  signed [7:0] mul_ln1352_16_fu_2422_p2;
wire   [3:0] mul_ln1352_17_fu_2435_p0;
wire  signed [7:0] mul_ln1352_17_fu_2435_p2;
wire   [3:0] mul_ln1352_18_fu_2448_p0;
wire  signed [7:0] mul_ln1352_18_fu_2448_p2;
wire   [3:0] mul_ln1352_19_fu_2461_p0;
wire  signed [7:0] mul_ln1352_19_fu_2461_p2;
wire   [3:0] mul_ln1352_20_fu_2474_p0;
wire  signed [7:0] mul_ln1352_20_fu_2474_p2;
wire   [3:0] mul_ln1352_21_fu_2487_p0;
wire   [3:0] mul_ln1352_22_fu_2496_p0;
wire  signed [7:0] mul_ln1352_22_fu_2496_p2;
wire   [3:0] mul_ln1352_23_fu_2509_p0;
wire  signed [7:0] mul_ln1352_23_fu_2509_p2;
wire  signed [8:0] sext_ln170_16_fu_2480_p1;
wire  signed [8:0] sext_ln170_17_fu_2502_p1;
wire  signed [8:0] sext_ln170_12_fu_2428_p1;
wire  signed [8:0] sext_ln170_15_fu_2467_p1;
wire  signed [8:0] sext_ln700_15_fu_2515_p1;
wire  signed [8:0] sext_ln170_13_fu_2441_p1;
wire   [8:0] add_ln700_20_fu_2531_p2;
wire  signed [9:0] sext_ln170_14_fu_2454_p1;
wire  signed [9:0] sext_ln700_18_fu_2537_p1;
wire   [3:0] mul_ln1352_24_fu_2550_p0;
wire  signed [7:0] mul_ln1352_24_fu_2550_p2;
wire   [3:0] mul_ln1352_25_fu_2563_p0;
wire  signed [7:0] mul_ln1352_25_fu_2563_p2;
wire   [3:0] mul_ln1352_26_fu_2576_p0;
wire  signed [7:0] mul_ln1352_26_fu_2576_p2;
wire   [3:0] mul_ln1352_27_fu_2589_p0;
wire  signed [7:0] mul_ln1352_27_fu_2589_p2;
wire   [3:0] mul_ln1352_28_fu_2602_p0;
wire  signed [7:0] mul_ln1352_28_fu_2602_p2;
wire   [3:0] mul_ln1352_29_fu_2615_p0;
wire   [3:0] mul_ln1352_30_fu_2624_p0;
wire  signed [7:0] mul_ln1352_30_fu_2624_p2;
wire   [3:0] mul_ln1352_31_fu_2637_p0;
wire  signed [7:0] mul_ln1352_31_fu_2637_p2;
wire  signed [8:0] sext_ln170_22_fu_2608_p1;
wire  signed [8:0] sext_ln170_23_fu_2630_p1;
wire  signed [8:0] sext_ln170_18_fu_2556_p1;
wire  signed [8:0] sext_ln170_21_fu_2595_p1;
wire  signed [8:0] sext_ln700_22_fu_2643_p1;
wire  signed [8:0] sext_ln170_19_fu_2569_p1;
wire   [8:0] add_ln700_28_fu_2659_p2;
wire  signed [9:0] sext_ln170_20_fu_2582_p1;
wire  signed [9:0] sext_ln700_25_fu_2665_p1;
wire   [31:0] nf_fu_2738_p2;
wire   [0:0] icmp_ln301_fu_2744_p2;
wire  signed [15:0] sext_ln700_fu_2803_p1;
wire   [15:0] select_ln271_3_fu_2796_p3;
wire   [15:0] add_ln700_fu_2806_p2;
wire  signed [15:0] sext_ln700_2_fu_2812_p1;
wire  signed [10:0] sext_ln700_3_fu_2821_p1;
wire  signed [10:0] sext_ln700_5_fu_2824_p1;
wire   [10:0] add_ln700_6_fu_2827_p2;
wire   [15:0] add_ln700_2_fu_2815_p2;
wire  signed [15:0] sext_ln700_6_fu_2833_p1;
wire  signed [15:0] sext_ln700_7_fu_2843_p1;
wire   [15:0] select_ln271_2_fu_2789_p3;
wire   [15:0] add_ln700_8_fu_2846_p2;
wire  signed [15:0] sext_ln700_9_fu_2852_p1;
wire  signed [10:0] sext_ln700_10_fu_2861_p1;
wire  signed [10:0] sext_ln700_12_fu_2864_p1;
wire   [10:0] add_ln700_14_fu_2867_p2;
wire   [15:0] add_ln700_10_fu_2855_p2;
wire  signed [15:0] sext_ln700_13_fu_2873_p1;
wire  signed [15:0] sext_ln700_14_fu_2883_p1;
wire   [15:0] select_ln271_1_fu_2782_p3;
wire   [15:0] add_ln700_16_fu_2886_p2;
wire  signed [15:0] sext_ln700_16_fu_2892_p1;
wire  signed [10:0] sext_ln700_17_fu_2901_p1;
wire  signed [10:0] sext_ln700_19_fu_2904_p1;
wire   [10:0] add_ln700_22_fu_2907_p2;
wire   [15:0] add_ln700_18_fu_2895_p2;
wire  signed [15:0] sext_ln700_20_fu_2913_p1;
wire  signed [15:0] sext_ln700_21_fu_2923_p1;
wire   [15:0] select_ln271_fu_2775_p3;
wire   [15:0] add_ln700_24_fu_2926_p2;
wire  signed [15:0] sext_ln700_23_fu_2932_p1;
wire  signed [10:0] sext_ln700_24_fu_2941_p1;
wire  signed [10:0] sext_ln700_26_fu_2944_p1;
wire   [10:0] add_ln700_30_fu_2947_p2;
wire   [15:0] add_ln700_26_fu_2935_p2;
wire  signed [15:0] sext_ln700_27_fu_2953_p1;
wire  signed [15:0] sext_ln142_fu_2983_p1;
wire  signed [15:0] sext_ln142_1_fu_2993_p1;
wire  signed [15:0] sext_ln142_2_fu_3099_p1;
wire  signed [15:0] sext_ln142_3_fu_3109_p1;
wire  signed [15:0] sext_ln142_4_fu_3119_p1;
wire  signed [15:0] sext_ln142_5_fu_3129_p1;
wire  signed [15:0] sext_ln142_6_fu_3139_p1;
wire  signed [15:0] sext_ln142_7_fu_3149_p1;
wire  signed [15:0] sext_ln142_8_fu_3159_p1;
wire  signed [15:0] sext_ln142_9_fu_3169_p1;
wire  signed [15:0] sext_ln142_10_fu_3179_p1;
wire  signed [15:0] sext_ln142_11_fu_3189_p1;
wire   [0:0] xor_ln899_3_fu_3367_p2;
wire   [0:0] xor_ln899_4_fu_3376_p2;
wire   [0:0] xor_ln899_5_fu_3385_p2;
wire   [0:0] xor_ln899_6_fu_3394_p2;
wire   [0:0] xor_ln899_7_fu_3403_p2;
wire   [0:0] xor_ln899_8_fu_3412_p2;
wire   [0:0] xor_ln899_9_fu_3421_p2;
wire   [0:0] xor_ln899_10_fu_3430_p2;
wire   [0:0] xor_ln899_11_fu_3439_p2;
wire   [0:0] xor_ln899_12_fu_3448_p2;
wire   [0:0] xor_ln899_13_fu_3457_p2;
wire   [1:0] zext_ln142_3_fu_3372_p1;
wire   [1:0] zext_ln142_4_fu_3381_p1;
wire   [1:0] add_ln700_34_fu_3466_p2;
wire   [1:0] zext_ln142_5_fu_3390_p1;
wire   [1:0] zext_ln142_6_fu_3399_p1;
wire   [1:0] add_ln700_35_fu_3476_p2;
wire   [2:0] zext_ln700_3_fu_3482_p1;
wire   [2:0] zext_ln700_2_fu_3472_p1;
wire   [1:0] zext_ln142_8_fu_3417_p1;
wire   [1:0] zext_ln142_9_fu_3426_p1;
wire   [1:0] add_ln700_38_fu_3492_p2;
wire   [1:0] zext_ln142_7_fu_3408_p1;
wire   [1:0] add_ln700_39_fu_3498_p2;
wire   [1:0] zext_ln142_10_fu_3435_p1;
wire   [1:0] zext_ln142_11_fu_3444_p1;
wire   [1:0] add_ln700_40_fu_3508_p2;
wire   [1:0] zext_ln142_12_fu_3453_p1;
wire   [1:0] zext_ln700_fu_3462_p1;
wire   [1:0] add_ln700_41_fu_3518_p2;
wire   [2:0] zext_ln700_7_fu_3524_p1;
wire   [2:0] zext_ln700_6_fu_3514_p1;
wire   [2:0] add_ln700_42_fu_3528_p2;
wire   [2:0] zext_ln700_5_fu_3504_p1;
wire   [0:0] xor_ln899_17_fu_3540_p2;
wire   [0:0] xor_ln899_18_fu_3549_p2;
wire   [0:0] xor_ln899_19_fu_3558_p2;
wire   [0:0] xor_ln899_20_fu_3567_p2;
wire   [0:0] xor_ln899_21_fu_3576_p2;
wire   [0:0] xor_ln899_22_fu_3585_p2;
wire   [0:0] xor_ln899_23_fu_3594_p2;
wire   [0:0] xor_ln899_24_fu_3603_p2;
wire   [0:0] xor_ln899_25_fu_3612_p2;
wire   [0:0] xor_ln899_26_fu_3621_p2;
wire   [0:0] xor_ln899_27_fu_3630_p2;
wire   [1:0] zext_ln142_15_fu_3545_p1;
wire   [1:0] zext_ln142_16_fu_3554_p1;
wire   [1:0] add_ln700_47_fu_3639_p2;
wire   [1:0] zext_ln142_17_fu_3563_p1;
wire   [1:0] zext_ln142_18_fu_3572_p1;
wire   [1:0] add_ln700_48_fu_3649_p2;
wire   [2:0] zext_ln700_12_fu_3655_p1;
wire   [2:0] zext_ln700_11_fu_3645_p1;
wire   [1:0] zext_ln142_20_fu_3590_p1;
wire   [1:0] zext_ln142_21_fu_3599_p1;
wire   [1:0] add_ln700_51_fu_3665_p2;
wire   [1:0] zext_ln142_19_fu_3581_p1;
wire   [1:0] add_ln700_52_fu_3671_p2;
wire   [1:0] zext_ln142_22_fu_3608_p1;
wire   [1:0] zext_ln142_23_fu_3617_p1;
wire   [1:0] add_ln700_53_fu_3681_p2;
wire   [1:0] zext_ln142_24_fu_3626_p1;
wire   [1:0] zext_ln700_9_fu_3635_p1;
wire   [1:0] add_ln700_54_fu_3691_p2;
wire   [2:0] zext_ln700_16_fu_3697_p1;
wire   [2:0] zext_ln700_15_fu_3687_p1;
wire   [2:0] add_ln700_55_fu_3701_p2;
wire   [2:0] zext_ln700_14_fu_3677_p1;
wire   [0:0] xor_ln899_31_fu_3713_p2;
wire   [0:0] xor_ln899_32_fu_3722_p2;
wire   [0:0] xor_ln899_33_fu_3731_p2;
wire   [0:0] xor_ln899_34_fu_3740_p2;
wire   [0:0] xor_ln899_35_fu_3749_p2;
wire   [0:0] xor_ln899_36_fu_3758_p2;
wire   [0:0] xor_ln899_37_fu_3767_p2;
wire   [0:0] xor_ln899_38_fu_3776_p2;
wire   [0:0] xor_ln899_39_fu_3785_p2;
wire   [0:0] xor_ln899_40_fu_3794_p2;
wire   [0:0] xor_ln899_41_fu_3803_p2;
wire   [1:0] zext_ln142_27_fu_3718_p1;
wire   [1:0] zext_ln142_28_fu_3727_p1;
wire   [1:0] add_ln700_60_fu_3812_p2;
wire   [1:0] zext_ln142_29_fu_3736_p1;
wire   [1:0] zext_ln142_30_fu_3745_p1;
wire   [1:0] add_ln700_61_fu_3822_p2;
wire   [2:0] zext_ln700_21_fu_3828_p1;
wire   [2:0] zext_ln700_20_fu_3818_p1;
wire   [1:0] zext_ln142_32_fu_3763_p1;
wire   [1:0] zext_ln142_33_fu_3772_p1;
wire   [1:0] add_ln700_64_fu_3838_p2;
wire   [1:0] zext_ln142_31_fu_3754_p1;
wire   [1:0] add_ln700_65_fu_3844_p2;
wire   [1:0] zext_ln142_34_fu_3781_p1;
wire   [1:0] zext_ln142_35_fu_3790_p1;
wire   [1:0] add_ln700_66_fu_3854_p2;
wire   [1:0] zext_ln142_36_fu_3799_p1;
wire   [1:0] zext_ln700_18_fu_3808_p1;
wire   [1:0] add_ln700_67_fu_3864_p2;
wire   [2:0] zext_ln700_25_fu_3870_p1;
wire   [2:0] zext_ln700_24_fu_3860_p1;
wire   [2:0] add_ln700_68_fu_3874_p2;
wire   [2:0] zext_ln700_23_fu_3850_p1;
wire   [0:0] xor_ln899_45_fu_3886_p2;
wire   [0:0] xor_ln899_46_fu_3895_p2;
wire   [0:0] xor_ln899_47_fu_3904_p2;
wire   [0:0] xor_ln899_48_fu_3913_p2;
wire   [0:0] xor_ln899_49_fu_3922_p2;
wire   [0:0] xor_ln899_50_fu_3931_p2;
wire   [0:0] xor_ln899_51_fu_3940_p2;
wire   [0:0] xor_ln899_52_fu_3949_p2;
wire   [0:0] xor_ln899_53_fu_3958_p2;
wire   [0:0] xor_ln899_54_fu_3967_p2;
wire   [0:0] xor_ln899_55_fu_3976_p2;
wire   [1:0] zext_ln142_39_fu_3891_p1;
wire   [1:0] zext_ln142_40_fu_3900_p1;
wire   [1:0] add_ln700_73_fu_3985_p2;
wire   [1:0] zext_ln142_41_fu_3909_p1;
wire   [1:0] zext_ln142_42_fu_3918_p1;
wire   [1:0] add_ln700_74_fu_3995_p2;
wire   [2:0] zext_ln700_30_fu_4001_p1;
wire   [2:0] zext_ln700_29_fu_3991_p1;
wire   [1:0] zext_ln142_44_fu_3936_p1;
wire   [1:0] zext_ln142_45_fu_3945_p1;
wire   [1:0] add_ln700_77_fu_4011_p2;
wire   [1:0] zext_ln142_43_fu_3927_p1;
wire   [1:0] add_ln700_78_fu_4017_p2;
wire   [1:0] zext_ln142_46_fu_3954_p1;
wire   [1:0] zext_ln142_47_fu_3963_p1;
wire   [1:0] add_ln700_79_fu_4027_p2;
wire   [1:0] zext_ln142_48_fu_3972_p1;
wire   [1:0] zext_ln700_27_fu_3981_p1;
wire   [1:0] add_ln700_80_fu_4037_p2;
wire   [2:0] zext_ln700_34_fu_4043_p1;
wire   [2:0] zext_ln700_33_fu_4033_p1;
wire   [2:0] add_ln700_81_fu_4047_p2;
wire   [2:0] zext_ln700_32_fu_4023_p1;
wire   [0:0] xor_ln899_fu_4059_p2;
wire   [0:0] xor_ln899_1_fu_4072_p2;
wire   [0:0] xor_ln899_2_fu_4081_p2;
wire   [1:0] zext_ln142_1_fu_4077_p1;
wire   [1:0] zext_ln142_2_fu_4086_p1;
wire   [1:0] add_ln700_32_fu_4090_p2;
wire   [3:0] zext_ln700_1_fu_4096_p1;
wire   [3:0] select_ln700_fu_4064_p3;
wire   [3:0] zext_ln700_4_fu_4106_p1;
wire   [3:0] add_ln700_33_fu_4100_p2;
wire   [3:0] zext_ln700_8_fu_4115_p1;
wire   [3:0] add_ln700_37_fu_4109_p2;
wire   [0:0] xor_ln899_14_fu_4124_p2;
wire   [0:0] xor_ln899_15_fu_4137_p2;
wire   [0:0] xor_ln899_16_fu_4146_p2;
wire   [1:0] zext_ln142_13_fu_4142_p1;
wire   [1:0] zext_ln142_14_fu_4151_p1;
wire   [1:0] add_ln700_45_fu_4155_p2;
wire   [3:0] zext_ln700_10_fu_4161_p1;
wire   [3:0] select_ln700_1_fu_4129_p3;
wire   [3:0] zext_ln700_13_fu_4171_p1;
wire   [3:0] add_ln700_46_fu_4165_p2;
wire   [3:0] zext_ln700_17_fu_4180_p1;
wire   [3:0] add_ln700_50_fu_4174_p2;
wire   [0:0] xor_ln899_28_fu_4189_p2;
wire   [0:0] xor_ln899_29_fu_4202_p2;
wire   [0:0] xor_ln899_30_fu_4211_p2;
wire   [1:0] zext_ln142_25_fu_4207_p1;
wire   [1:0] zext_ln142_26_fu_4216_p1;
wire   [1:0] add_ln700_58_fu_4220_p2;
wire   [3:0] zext_ln700_19_fu_4226_p1;
wire   [3:0] select_ln700_2_fu_4194_p3;
wire   [3:0] zext_ln700_22_fu_4236_p1;
wire   [3:0] add_ln700_59_fu_4230_p2;
wire   [3:0] zext_ln700_26_fu_4245_p1;
wire   [3:0] add_ln700_63_fu_4239_p2;
wire   [0:0] xor_ln899_42_fu_4254_p2;
wire   [0:0] xor_ln899_43_fu_4267_p2;
wire   [0:0] xor_ln899_44_fu_4276_p2;
wire   [1:0] zext_ln142_37_fu_4272_p1;
wire   [1:0] zext_ln142_38_fu_4281_p1;
wire   [1:0] add_ln700_71_fu_4285_p2;
wire   [3:0] zext_ln700_28_fu_4291_p1;
wire   [3:0] select_ln700_3_fu_4259_p3;
wire   [3:0] zext_ln700_31_fu_4301_p1;
wire   [3:0] add_ln700_72_fu_4295_p2;
wire   [3:0] zext_ln700_35_fu_4310_p1;
wire   [3:0] add_ln700_76_fu_4304_p2;
wire   [3:0] add_ln700_83_fu_4313_p2;
wire   [3:0] add_ln700_70_fu_4248_p2;
wire   [3:0] add_ln700_57_fu_4183_p2;
wire   [3:0] add_ln700_44_fu_4118_p2;
wire    ap_CS_fsm_state7;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
end

StreamingFCLayer_Batch_3_Matrix_Vector_Actbkb #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_55_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_55_address0),
    .ce0(threshs_m_thresholds_55_ce0),
    .q0(threshs_m_thresholds_55_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actcud #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_54_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_54_address0),
    .ce0(threshs_m_thresholds_54_ce0),
    .q0(threshs_m_thresholds_54_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActdEe #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_49_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_49_address0),
    .ce0(threshs_m_thresholds_49_ce0),
    .q0(threshs_m_thresholds_49_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActeOg #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_48_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_48_address0),
    .ce0(threshs_m_thresholds_48_ce0),
    .q0(threshs_m_thresholds_48_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActfYi #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_47_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_47_address0),
    .ce0(threshs_m_thresholds_47_ce0),
    .q0(threshs_m_thresholds_47_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actg8j #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_46_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_46_address0),
    .ce0(threshs_m_thresholds_46_ce0),
    .q0(threshs_m_thresholds_46_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Acthbi #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_45_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_45_address0),
    .ce0(threshs_m_thresholds_45_ce0),
    .q0(threshs_m_thresholds_45_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actibs #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_44_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_44_address0),
    .ce0(threshs_m_thresholds_44_ce0),
    .q0(threshs_m_thresholds_44_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActjbC #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_43_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_43_address0),
    .ce0(threshs_m_thresholds_43_ce0),
    .q0(threshs_m_thresholds_43_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActkbM #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_42_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_42_address0),
    .ce0(threshs_m_thresholds_42_ce0),
    .q0(threshs_m_thresholds_42_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActlbW #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_53_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_53_address0),
    .ce0(threshs_m_thresholds_53_ce0),
    .q0(threshs_m_thresholds_53_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actmb6 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_52_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_52_address0),
    .ce0(threshs_m_thresholds_52_ce0),
    .q0(threshs_m_thresholds_52_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actncg #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_51_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_51_address0),
    .ce0(threshs_m_thresholds_51_ce0),
    .q0(threshs_m_thresholds_51_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actocq #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_50_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_50_address0),
    .ce0(threshs_m_thresholds_50_ce0),
    .q0(threshs_m_thresholds_50_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActpcA #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_41_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_41_address0),
    .ce0(threshs_m_thresholds_41_ce0),
    .q0(threshs_m_thresholds_41_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActqcK #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_40_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_40_address0),
    .ce0(threshs_m_thresholds_40_ce0),
    .q0(threshs_m_thresholds_40_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActrcU #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_35_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_35_address0),
    .ce0(threshs_m_thresholds_35_ce0),
    .q0(threshs_m_thresholds_35_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actsc4 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_34_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_34_address0),
    .ce0(threshs_m_thresholds_34_ce0),
    .q0(threshs_m_thresholds_34_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Acttde #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_33_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_33_address0),
    .ce0(threshs_m_thresholds_33_ce0),
    .q0(threshs_m_thresholds_33_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actudo #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_32_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_32_address0),
    .ce0(threshs_m_thresholds_32_ce0),
    .q0(threshs_m_thresholds_32_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actvdy #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_31_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_31_address0),
    .ce0(threshs_m_thresholds_31_ce0),
    .q0(threshs_m_thresholds_31_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActwdI #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_30_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_30_address0),
    .ce0(threshs_m_thresholds_30_ce0),
    .q0(threshs_m_thresholds_30_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActxdS #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_29_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_29_address0),
    .ce0(threshs_m_thresholds_29_ce0),
    .q0(threshs_m_thresholds_29_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actyd2 #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_28_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_28_address0),
    .ce0(threshs_m_thresholds_28_ce0),
    .q0(threshs_m_thresholds_28_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Actzec #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_39_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_39_address0),
    .ce0(threshs_m_thresholds_39_ce0),
    .q0(threshs_m_thresholds_39_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActAem #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_38_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_38_address0),
    .ce0(threshs_m_thresholds_38_ce0),
    .q0(threshs_m_thresholds_38_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActBew #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_37_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_37_address0),
    .ce0(threshs_m_thresholds_37_ce0),
    .q0(threshs_m_thresholds_37_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActCeG #(
    .DataWidth( 15 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_36_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_36_address0),
    .ce0(threshs_m_thresholds_36_ce0),
    .q0(threshs_m_thresholds_36_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActDeQ #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_27_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_27_address0),
    .ce0(threshs_m_thresholds_27_ce0),
    .q0(threshs_m_thresholds_27_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActEe0 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_26_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_26_address0),
    .ce0(threshs_m_thresholds_26_ce0),
    .q0(threshs_m_thresholds_26_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActFfa #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_21_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_21_address0),
    .ce0(threshs_m_thresholds_21_ce0),
    .q0(threshs_m_thresholds_21_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActGfk #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_20_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_20_address0),
    .ce0(threshs_m_thresholds_20_ce0),
    .q0(threshs_m_thresholds_20_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActHfu #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_19_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_19_address0),
    .ce0(threshs_m_thresholds_19_ce0),
    .q0(threshs_m_thresholds_19_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActIfE #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_18_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_18_address0),
    .ce0(threshs_m_thresholds_18_ce0),
    .q0(threshs_m_thresholds_18_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActJfO #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_17_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_17_address0),
    .ce0(threshs_m_thresholds_17_ce0),
    .q0(threshs_m_thresholds_17_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActKfY #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_16_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_16_address0),
    .ce0(threshs_m_thresholds_16_ce0),
    .q0(threshs_m_thresholds_16_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActLf8 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_15_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_15_address0),
    .ce0(threshs_m_thresholds_15_ce0),
    .q0(threshs_m_thresholds_15_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActMgi #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_14_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_14_address0),
    .ce0(threshs_m_thresholds_14_ce0),
    .q0(threshs_m_thresholds_14_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActNgs #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_25_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_25_address0),
    .ce0(threshs_m_thresholds_25_ce0),
    .q0(threshs_m_thresholds_25_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActOgC #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_24_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_24_address0),
    .ce0(threshs_m_thresholds_24_ce0),
    .q0(threshs_m_thresholds_24_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActPgM #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_23_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_23_address0),
    .ce0(threshs_m_thresholds_23_ce0),
    .q0(threshs_m_thresholds_23_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActQgW #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_22_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_22_address0),
    .ce0(threshs_m_thresholds_22_ce0),
    .q0(threshs_m_thresholds_22_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActRg6 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_13_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_13_address0),
    .ce0(threshs_m_thresholds_13_ce0),
    .q0(threshs_m_thresholds_13_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActShg #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_12_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_12_address0),
    .ce0(threshs_m_thresholds_12_ce0),
    .q0(threshs_m_thresholds_12_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActThq #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_7_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_7_address0),
    .ce0(threshs_m_thresholds_7_ce0),
    .q0(threshs_m_thresholds_7_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActUhA #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_6_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_6_address0),
    .ce0(threshs_m_thresholds_6_ce0),
    .q0(threshs_m_thresholds_6_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActVhK #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_5_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_5_address0),
    .ce0(threshs_m_thresholds_5_ce0),
    .q0(threshs_m_thresholds_5_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActWhU #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_4_address0),
    .ce0(threshs_m_thresholds_4_ce0),
    .q0(threshs_m_thresholds_4_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActXh4 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_3_address0),
    .ce0(threshs_m_thresholds_3_ce0),
    .q0(threshs_m_thresholds_3_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActYie #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_2_address0),
    .ce0(threshs_m_thresholds_2_ce0),
    .q0(threshs_m_thresholds_2_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_ActZio #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_1_address0),
    .ce0(threshs_m_thresholds_1_ce0),
    .q0(threshs_m_thresholds_1_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Act0iy #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_address0),
    .ce0(threshs_m_thresholds_ce0),
    .q0(threshs_m_thresholds_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Act1iI #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_11_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_11_address0),
    .ce0(threshs_m_thresholds_11_ce0),
    .q0(threshs_m_thresholds_11_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Act2iS #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_10_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_10_address0),
    .ce0(threshs_m_thresholds_10_ce0),
    .q0(threshs_m_thresholds_10_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Act3i2 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_9_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_9_address0),
    .ce0(threshs_m_thresholds_9_ce0),
    .q0(threshs_m_thresholds_9_q0)
);

StreamingFCLayer_Batch_3_Matrix_Vector_Act4jc #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_8_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_8_address0),
    .ce0(threshs_m_thresholds_8_ce0),
    .q0(threshs_m_thresholds_8_q0)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_5jm #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 32 ),
    .din5_WIDTH( 32 ),
    .din6_WIDTH( 32 ),
    .din7_WIDTH( 32 ),
    .din8_WIDTH( 32 ),
    .din9_WIDTH( 32 ),
    .din10_WIDTH( 32 ),
    .din11_WIDTH( 32 ),
    .din12_WIDTH( 32 ),
    .din13_WIDTH( 32 ),
    .din14_WIDTH( 32 ),
    .din15_WIDTH( 32 ),
    .din16_WIDTH( 32 ),
    .din17_WIDTH( 32 ),
    .din18_WIDTH( 32 ),
    .din19_WIDTH( 32 ),
    .din20_WIDTH( 32 ),
    .din21_WIDTH( 32 ),
    .din22_WIDTH( 32 ),
    .din23_WIDTH( 32 ),
    .din24_WIDTH( 32 ),
    .din25_WIDTH( 32 ),
    .din26_WIDTH( 32 ),
    .din27_WIDTH( 32 ),
    .din28_WIDTH( 32 ),
    .din29_WIDTH( 32 ),
    .din30_WIDTH( 32 ),
    .din31_WIDTH( 32 ),
    .din32_WIDTH( 5 ),
    .dout_WIDTH( 32 ))
StreamingFCLayer_5jm_U1(
    .din0(tmp_V_fu_388),
    .din1(tmp_V_1_fu_392),
    .din2(tmp_V_2_fu_396),
    .din3(tmp_V_4_fu_400),
    .din4(tmp_V_5_fu_404),
    .din5(tmp_V_6_fu_408),
    .din6(tmp_V_7_fu_412),
    .din7(tmp_V_8_fu_416),
    .din8(tmp_V_9_fu_420),
    .din9(tmp_V_10_fu_424),
    .din10(tmp_V_11_fu_428),
    .din11(tmp_V_12_fu_432),
    .din12(tmp_V_13_fu_436),
    .din13(tmp_V_14_fu_440),
    .din14(tmp_V_15_fu_444),
    .din15(tmp_V_16_fu_448),
    .din16(tmp_V_17_fu_452),
    .din17(tmp_V_18_fu_456),
    .din18(tmp_V_19_fu_460),
    .din19(tmp_V_20_fu_464),
    .din20(tmp_V_21_fu_468),
    .din21(tmp_V_22_fu_472),
    .din22(tmp_V_23_fu_476),
    .din23(tmp_V_24_fu_480),
    .din24(tmp_V_25_fu_484),
    .din25(tmp_V_26_fu_488),
    .din26(tmp_V_27_fu_492),
    .din27(tmp_V_28_fu_496),
    .din28(tmp_V_29_fu_500),
    .din29(tmp_V_30_fu_504),
    .din30(tmp_V_31_fu_508),
    .din31(tmp_V_32_fu_512),
    .din32(inElem_V_1_fu_1483_p33),
    .dout(inElem_V_1_fu_1483_p34)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U2(
    .din0(mul_ln1352_fu_2068_p0),
    .din1(wgt_M_instance_0_V_reg_4630),
    .dout(mul_ln1352_fu_2068_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U3(
    .din0(mul_ln1352_1_fu_2095_p0),
    .din1(wgt_M_instance_1_V_reg_4635),
    .dout(mul_ln1352_1_fu_2095_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U4(
    .din0(mul_ln1352_2_fu_2122_p0),
    .din1(wgt_M_instance_2_V_reg_4640),
    .dout(mul_ln1352_2_fu_2122_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U5(
    .din0(mul_ln1352_3_fu_2149_p0),
    .din1(wgt_M_instance_3_V_reg_4645),
    .dout(mul_ln1352_3_fu_2149_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U6(
    .din0(mul_ln1352_4_fu_2176_p0),
    .din1(wgt_M_instance_4_V_reg_4650),
    .dout(mul_ln1352_4_fu_2176_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U7(
    .din0(mul_ln1352_5_fu_2203_p0),
    .din1(wgt_M_instance_5_V_reg_4655),
    .dout(mul_ln1352_5_fu_2203_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U8(
    .din0(mul_ln1352_6_fu_2226_p0),
    .din1(wgt_M_instance_6_V_reg_4660),
    .dout(mul_ln1352_6_fu_2226_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U9(
    .din0(mul_ln1352_7_fu_2253_p0),
    .din1(wgt_M_instance_7_V_reg_4665),
    .dout(mul_ln1352_7_fu_2253_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U10(
    .din0(mul_ln1352_8_fu_2294_p0),
    .din1(wgt_M_instance_0_V_1_reg_4670),
    .dout(mul_ln1352_8_fu_2294_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U11(
    .din0(mul_ln1352_9_fu_2307_p0),
    .din1(wgt_M_instance_1_V_1_reg_4675),
    .dout(mul_ln1352_9_fu_2307_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U12(
    .din0(mul_ln1352_10_fu_2320_p0),
    .din1(wgt_M_instance_2_V_1_reg_4680),
    .dout(mul_ln1352_10_fu_2320_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U13(
    .din0(mul_ln1352_11_fu_2333_p0),
    .din1(wgt_M_instance_3_V_1_reg_4685),
    .dout(mul_ln1352_11_fu_2333_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U14(
    .din0(mul_ln1352_12_fu_2346_p0),
    .din1(wgt_M_instance_4_V_1_reg_4690),
    .dout(mul_ln1352_12_fu_2346_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U15(
    .din0(mul_ln1352_13_fu_2359_p0),
    .din1(wgt_M_instance_5_V_1_reg_4695),
    .dout(mul_ln1352_13_fu_2359_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U16(
    .din0(mul_ln1352_14_fu_2368_p0),
    .din1(wgt_M_instance_6_V_1_reg_4700),
    .dout(mul_ln1352_14_fu_2368_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U17(
    .din0(mul_ln1352_15_fu_2381_p0),
    .din1(wgt_M_instance_7_V_1_reg_4705),
    .dout(mul_ln1352_15_fu_2381_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U18(
    .din0(mul_ln1352_16_fu_2422_p0),
    .din1(wgt_M_instance_0_V_2_reg_4710),
    .dout(mul_ln1352_16_fu_2422_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U19(
    .din0(mul_ln1352_17_fu_2435_p0),
    .din1(wgt_M_instance_1_V_2_reg_4715),
    .dout(mul_ln1352_17_fu_2435_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U20(
    .din0(mul_ln1352_18_fu_2448_p0),
    .din1(wgt_M_instance_2_V_2_reg_4720),
    .dout(mul_ln1352_18_fu_2448_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U21(
    .din0(mul_ln1352_19_fu_2461_p0),
    .din1(wgt_M_instance_3_V_2_reg_4725),
    .dout(mul_ln1352_19_fu_2461_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U22(
    .din0(mul_ln1352_20_fu_2474_p0),
    .din1(wgt_M_instance_4_V_2_reg_4730),
    .dout(mul_ln1352_20_fu_2474_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U23(
    .din0(mul_ln1352_21_fu_2487_p0),
    .din1(wgt_M_instance_5_V_2_reg_4735),
    .dout(mul_ln1352_21_fu_2487_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U24(
    .din0(mul_ln1352_22_fu_2496_p0),
    .din1(wgt_M_instance_6_V_2_reg_4740),
    .dout(mul_ln1352_22_fu_2496_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U25(
    .din0(mul_ln1352_23_fu_2509_p0),
    .din1(wgt_M_instance_7_V_2_reg_4745),
    .dout(mul_ln1352_23_fu_2509_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U26(
    .din0(mul_ln1352_24_fu_2550_p0),
    .din1(wgt_M_instance_0_V_3_reg_4750),
    .dout(mul_ln1352_24_fu_2550_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U27(
    .din0(mul_ln1352_25_fu_2563_p0),
    .din1(wgt_M_instance_1_V_3_reg_4755),
    .dout(mul_ln1352_25_fu_2563_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U28(
    .din0(mul_ln1352_26_fu_2576_p0),
    .din1(wgt_M_instance_2_V_3_reg_4760),
    .dout(mul_ln1352_26_fu_2576_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U29(
    .din0(mul_ln1352_27_fu_2589_p0),
    .din1(wgt_M_instance_3_V_3_reg_4765),
    .dout(mul_ln1352_27_fu_2589_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U30(
    .din0(mul_ln1352_28_fu_2602_p0),
    .din1(wgt_M_instance_4_V_3_reg_4770),
    .dout(mul_ln1352_28_fu_2602_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U31(
    .din0(mul_ln1352_29_fu_2615_p0),
    .din1(wgt_M_instance_5_V_3_reg_4775),
    .dout(mul_ln1352_29_fu_2615_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U32(
    .din0(mul_ln1352_30_fu_2624_p0),
    .din1(wgt_M_instance_6_V_3_reg_4780),
    .dout(mul_ln1352_30_fu_2624_p2)
);

StreamingFCLayer_Batch_3_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U33(
    .din0(mul_ln1352_31_fu_2637_p0),
    .din1(wgt_M_instance_7_V_3_reg_4785),
    .dout(mul_ln1352_31_fu_2637_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd0) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278 <= inElem_V_1_fu_1483_p34;
    end else if ((((trunc_ln321_fu_1553_p1 == 5'd14) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd15) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd16) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd17) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd18) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd19) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd20) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd21) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd22) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd23) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd24) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd25) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd26) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd27) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd28) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd29) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd30) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd31) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd2) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd3) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd4) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd5) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd6) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd7) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd8) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd9) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd10) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd11) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd12) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1553_p1 == 5'd13) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278 <= in_V_V_TDATA;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278 <= ap_phi_reg_pp0_iter0_act_m_val_V_reg_1278;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_reg_1267 <= i_fu_1365_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_reg_1267 <= 13'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_4790 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        nf_assign_fu_516 <= select_ln301_fu_2750_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        nf_assign_fu_516 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_2046_p2 == 1'd0) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        sf_1_fu_384 <= sf_fu_2040_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_2046_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        sf_1_fu_384 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        accu_V_0_0_0_fu_368 <= accu_0_0_V_fu_2837_p2;
        accu_V_0_1_0_fu_372 <= accu_0_1_V_fu_2877_p2;
        accu_V_0_2_0_fu_376 <= accu_0_2_V_fu_2917_p2;
        accu_V_0_3_0_fu_380 <= accu_0_3_V_fu_2957_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln700_11_reg_4824 <= add_ln700_11_fu_2397_p2;
        add_ln700_13_reg_4829 <= add_ln700_13_fu_2413_p2;
        add_ln700_17_reg_4839 <= add_ln700_17_fu_2519_p2;
        add_ln700_19_reg_4844 <= add_ln700_19_fu_2525_p2;
        add_ln700_1_reg_4799 <= add_ln700_1_fu_2263_p2;
        add_ln700_21_reg_4849 <= add_ln700_21_fu_2541_p2;
        add_ln700_25_reg_4859 <= add_ln700_25_fu_2647_p2;
        add_ln700_27_reg_4864 <= add_ln700_27_fu_2653_p2;
        add_ln700_29_reg_4869 <= add_ln700_29_fu_2669_p2;
        add_ln700_3_reg_4804 <= add_ln700_3_fu_2269_p2;
        add_ln700_5_reg_4809 <= add_ln700_5_fu_2285_p2;
        add_ln700_9_reg_4819 <= add_ln700_9_fu_2391_p2;
        icmp_ln271_reg_4622_pp0_iter1_reg <= icmp_ln271_reg_4622;
        icmp_ln289_reg_4790_pp0_iter1_reg <= icmp_ln289_reg_4790;
        mul_ln1352_13_reg_4814 <= mul_ln1352_13_fu_2359_p2;
        mul_ln1352_21_reg_4834 <= mul_ln1352_21_fu_2487_p2;
        mul_ln1352_29_reg_4854 <= mul_ln1352_29_fu_2615_p2;
        mul_ln1352_5_reg_4794 <= mul_ln1352_5_fu_2203_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_4790_pp0_iter2_reg == 1'd1))) begin
        add_ln700_36_reg_5434 <= add_ln700_36_fu_3486_p2;
        add_ln700_43_reg_5439 <= add_ln700_43_fu_3534_p2;
        add_ln700_49_reg_5444 <= add_ln700_49_fu_3659_p2;
        add_ln700_56_reg_5449 <= add_ln700_56_fu_3707_p2;
        add_ln700_62_reg_5454 <= add_ln700_62_fu_3832_p2;
        add_ln700_69_reg_5459 <= add_ln700_69_fu_3880_p2;
        add_ln700_75_reg_5464 <= add_ln700_75_fu_4005_p2;
        add_ln700_82_reg_5469 <= add_ln700_82_fu_4053_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_1359_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln271_reg_4622 <= icmp_ln271_fu_1720_p2;
        icmp_ln289_reg_4790 <= icmp_ln289_fu_2046_p2;
        wgt_M_instance_0_V_1_reg_4670 <= {{weight_V_V_TDATA[35:32]}};
        wgt_M_instance_0_V_2_reg_4710 <= {{weight_V_V_TDATA[67:64]}};
        wgt_M_instance_0_V_3_reg_4750 <= {{weight_V_V_TDATA[99:96]}};
        wgt_M_instance_0_V_reg_4630 <= wgt_M_instance_0_V_fu_1726_p1;
        wgt_M_instance_1_V_1_reg_4675 <= {{weight_V_V_TDATA[39:36]}};
        wgt_M_instance_1_V_2_reg_4715 <= {{weight_V_V_TDATA[71:68]}};
        wgt_M_instance_1_V_3_reg_4755 <= {{weight_V_V_TDATA[103:100]}};
        wgt_M_instance_1_V_reg_4635 <= {{weight_V_V_TDATA[7:4]}};
        wgt_M_instance_2_V_1_reg_4680 <= {{weight_V_V_TDATA[43:40]}};
        wgt_M_instance_2_V_2_reg_4720 <= {{weight_V_V_TDATA[75:72]}};
        wgt_M_instance_2_V_3_reg_4760 <= {{weight_V_V_TDATA[107:104]}};
        wgt_M_instance_2_V_reg_4640 <= {{weight_V_V_TDATA[11:8]}};
        wgt_M_instance_3_V_1_reg_4685 <= {{weight_V_V_TDATA[47:44]}};
        wgt_M_instance_3_V_2_reg_4725 <= {{weight_V_V_TDATA[79:76]}};
        wgt_M_instance_3_V_3_reg_4765 <= {{weight_V_V_TDATA[111:108]}};
        wgt_M_instance_3_V_reg_4645 <= {{weight_V_V_TDATA[15:12]}};
        wgt_M_instance_4_V_1_reg_4690 <= {{weight_V_V_TDATA[51:48]}};
        wgt_M_instance_4_V_2_reg_4730 <= {{weight_V_V_TDATA[83:80]}};
        wgt_M_instance_4_V_3_reg_4770 <= {{weight_V_V_TDATA[115:112]}};
        wgt_M_instance_4_V_reg_4650 <= {{weight_V_V_TDATA[19:16]}};
        wgt_M_instance_5_V_1_reg_4695 <= {{weight_V_V_TDATA[55:52]}};
        wgt_M_instance_5_V_2_reg_4735 <= {{weight_V_V_TDATA[87:84]}};
        wgt_M_instance_5_V_3_reg_4775 <= {{weight_V_V_TDATA[119:116]}};
        wgt_M_instance_5_V_reg_4655 <= {{weight_V_V_TDATA[23:20]}};
        wgt_M_instance_6_V_1_reg_4700 <= {{weight_V_V_TDATA[59:56]}};
        wgt_M_instance_6_V_2_reg_4740 <= {{weight_V_V_TDATA[91:88]}};
        wgt_M_instance_6_V_3_reg_4780 <= {{weight_V_V_TDATA[123:120]}};
        wgt_M_instance_6_V_reg_4660 <= {{weight_V_V_TDATA[27:24]}};
        wgt_M_instance_7_V_1_reg_4705 <= {{weight_V_V_TDATA[63:60]}};
        wgt_M_instance_7_V_2_reg_4745 <= {{weight_V_V_TDATA[95:92]}};
        wgt_M_instance_7_V_3_reg_4785 <= {{weight_V_V_TDATA[127:124]}};
        wgt_M_instance_7_V_reg_4665 <= {{weight_V_V_TDATA[31:28]}};
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln289_reg_4790_pp0_iter2_reg <= icmp_ln289_reg_4790_pp0_iter1_reg;
        icmp_ln289_reg_4790_pp0_iter3_reg <= icmp_ln289_reg_4790_pp0_iter2_reg;
        icmp_ln899_14_reg_5224_pp0_iter3_reg <= icmp_ln899_14_reg_5224;
        icmp_ln899_15_reg_5229_pp0_iter3_reg <= icmp_ln899_15_reg_5229;
        icmp_ln899_16_reg_5234_pp0_iter3_reg <= icmp_ln899_16_reg_5234;
        icmp_ln899_1_reg_5159_pp0_iter3_reg <= icmp_ln899_1_reg_5159;
        icmp_ln899_28_reg_5294_pp0_iter3_reg <= icmp_ln899_28_reg_5294;
        icmp_ln899_29_reg_5299_pp0_iter3_reg <= icmp_ln899_29_reg_5299;
        icmp_ln899_2_reg_5164_pp0_iter3_reg <= icmp_ln899_2_reg_5164;
        icmp_ln899_30_reg_5304_pp0_iter3_reg <= icmp_ln899_30_reg_5304;
        icmp_ln899_42_reg_5364_pp0_iter3_reg <= icmp_ln899_42_reg_5364;
        icmp_ln899_43_reg_5369_pp0_iter3_reg <= icmp_ln899_43_reg_5369;
        icmp_ln899_44_reg_5374_pp0_iter3_reg <= icmp_ln899_44_reg_5374;
        icmp_ln899_reg_5154_pp0_iter3_reg <= icmp_ln899_reg_5154;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_4790_pp0_iter1_reg == 1'd1))) begin
        icmp_ln899_10_reg_5204 <= icmp_ln899_10_fu_3051_p2;
        icmp_ln899_11_reg_5209 <= icmp_ln899_11_fu_3057_p2;
        icmp_ln899_12_reg_5214 <= icmp_ln899_12_fu_3063_p2;
        icmp_ln899_13_reg_5219 <= icmp_ln899_13_fu_3069_p2;
        icmp_ln899_14_reg_5224 <= icmp_ln899_14_fu_3075_p2;
        icmp_ln899_15_reg_5229 <= icmp_ln899_15_fu_3081_p2;
        icmp_ln899_16_reg_5234 <= icmp_ln899_16_fu_3087_p2;
        icmp_ln899_17_reg_5239 <= icmp_ln899_17_fu_3093_p2;
        icmp_ln899_18_reg_5244 <= icmp_ln899_18_fu_3103_p2;
        icmp_ln899_19_reg_5249 <= icmp_ln899_19_fu_3113_p2;
        icmp_ln899_1_reg_5159 <= icmp_ln899_1_fu_2997_p2;
        icmp_ln899_20_reg_5254 <= icmp_ln899_20_fu_3123_p2;
        icmp_ln899_21_reg_5259 <= icmp_ln899_21_fu_3133_p2;
        icmp_ln899_22_reg_5264 <= icmp_ln899_22_fu_3143_p2;
        icmp_ln899_23_reg_5269 <= icmp_ln899_23_fu_3153_p2;
        icmp_ln899_24_reg_5274 <= icmp_ln899_24_fu_3163_p2;
        icmp_ln899_25_reg_5279 <= icmp_ln899_25_fu_3173_p2;
        icmp_ln899_26_reg_5284 <= icmp_ln899_26_fu_3183_p2;
        icmp_ln899_27_reg_5289 <= icmp_ln899_27_fu_3193_p2;
        icmp_ln899_28_reg_5294 <= icmp_ln899_28_fu_3199_p2;
        icmp_ln899_29_reg_5299 <= icmp_ln899_29_fu_3205_p2;
        icmp_ln899_2_reg_5164 <= icmp_ln899_2_fu_3003_p2;
        icmp_ln899_30_reg_5304 <= icmp_ln899_30_fu_3211_p2;
        icmp_ln899_31_reg_5309 <= icmp_ln899_31_fu_3217_p2;
        icmp_ln899_32_reg_5314 <= icmp_ln899_32_fu_3223_p2;
        icmp_ln899_33_reg_5319 <= icmp_ln899_33_fu_3229_p2;
        icmp_ln899_34_reg_5324 <= icmp_ln899_34_fu_3235_p2;
        icmp_ln899_35_reg_5329 <= icmp_ln899_35_fu_3241_p2;
        icmp_ln899_36_reg_5334 <= icmp_ln899_36_fu_3247_p2;
        icmp_ln899_37_reg_5339 <= icmp_ln899_37_fu_3253_p2;
        icmp_ln899_38_reg_5344 <= icmp_ln899_38_fu_3259_p2;
        icmp_ln899_39_reg_5349 <= icmp_ln899_39_fu_3265_p2;
        icmp_ln899_3_reg_5169 <= icmp_ln899_3_fu_3009_p2;
        icmp_ln899_40_reg_5354 <= icmp_ln899_40_fu_3271_p2;
        icmp_ln899_41_reg_5359 <= icmp_ln899_41_fu_3277_p2;
        icmp_ln899_42_reg_5364 <= icmp_ln899_42_fu_3283_p2;
        icmp_ln899_43_reg_5369 <= icmp_ln899_43_fu_3289_p2;
        icmp_ln899_44_reg_5374 <= icmp_ln899_44_fu_3295_p2;
        icmp_ln899_45_reg_5379 <= icmp_ln899_45_fu_3301_p2;
        icmp_ln899_46_reg_5384 <= icmp_ln899_46_fu_3307_p2;
        icmp_ln899_47_reg_5389 <= icmp_ln899_47_fu_3313_p2;
        icmp_ln899_48_reg_5394 <= icmp_ln899_48_fu_3319_p2;
        icmp_ln899_49_reg_5399 <= icmp_ln899_49_fu_3325_p2;
        icmp_ln899_4_reg_5174 <= icmp_ln899_4_fu_3015_p2;
        icmp_ln899_50_reg_5404 <= icmp_ln899_50_fu_3331_p2;
        icmp_ln899_51_reg_5409 <= icmp_ln899_51_fu_3337_p2;
        icmp_ln899_52_reg_5414 <= icmp_ln899_52_fu_3343_p2;
        icmp_ln899_53_reg_5419 <= icmp_ln899_53_fu_3349_p2;
        icmp_ln899_54_reg_5424 <= icmp_ln899_54_fu_3355_p2;
        icmp_ln899_55_reg_5429 <= icmp_ln899_55_fu_3361_p2;
        icmp_ln899_5_reg_5179 <= icmp_ln899_5_fu_3021_p2;
        icmp_ln899_6_reg_5184 <= icmp_ln899_6_fu_3027_p2;
        icmp_ln899_7_reg_5189 <= icmp_ln899_7_fu_3033_p2;
        icmp_ln899_8_reg_5194 <= icmp_ln899_8_fu_3039_p2;
        icmp_ln899_9_reg_5199 <= icmp_ln899_9_fu_3045_p2;
        icmp_ln899_reg_5154 <= icmp_ln899_fu_2987_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd9) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_10_fu_424 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd10) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_11_fu_428 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd11) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_12_fu_432 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd12) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_13_fu_436 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd13) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_14_fu_440 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd14) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_15_fu_444 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd15) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_16_fu_448 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd16) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_17_fu_452 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd17) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_18_fu_456 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd18) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_19_fu_460 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_1_fu_392 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd19) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_20_fu_464 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd20) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_21_fu_468 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd21) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_22_fu_472 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd22) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_23_fu_476 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd23) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_24_fu_480 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd24) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_25_fu_484 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd25) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_26_fu_488 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd26) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_27_fu_492 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd27) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_28_fu_496 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd28) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_29_fu_500 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd2) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_2_fu_396 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd29) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_30_fu_504 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd30) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_31_fu_508 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd31) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_32_fu_512 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd3) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_4_fu_400 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd4) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_5_fu_404 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd5) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_6_fu_408 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd6) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_7_fu_412 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd7) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_8_fu_416 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd8) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_9_fu_420 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1553_p1 == 5'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_fu_388 <= in_V_V_TDATA;
    end
end

always @ (*) begin
    if ((icmp_ln248_fu_1359_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state7) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_4790 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_sig_allocacmp_nf_assign_load_1 = select_ln301_fu_2750_p3;
    end else begin
        ap_sig_allocacmp_nf_assign_load_1 = nf_assign_fu_516;
    end
end

always @ (*) begin
    if (((icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op98_read_state2 == 1'b1))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_4790_pp0_iter3_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_4790_pp0_iter3_reg == 1'd1) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_10_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_10_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_11_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_11_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_12_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_12_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_13_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_13_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_14_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_14_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_15_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_15_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_16_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_16_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_17_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_17_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_18_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_18_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_19_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_19_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_1_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_1_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_20_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_20_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_21_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_21_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_22_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_22_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_23_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_23_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_24_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_24_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_25_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_25_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_26_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_26_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_27_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_27_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_28_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_28_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_29_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_29_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_2_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_2_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_30_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_30_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_31_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_31_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_32_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_32_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_33_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_33_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_34_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_34_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_35_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_35_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_36_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_36_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_37_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_37_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_38_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_38_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_39_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_39_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_3_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_3_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_40_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_40_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_41_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_41_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_42_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_42_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_43_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_43_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_44_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_44_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_45_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_45_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_46_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_46_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_47_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_47_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_48_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_48_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_49_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_49_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_4_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_4_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_50_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_50_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_51_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_51_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_52_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_52_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_53_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_53_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_54_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_54_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_55_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_55_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_5_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_5_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_6_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_6_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_7_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_7_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_8_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_8_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_9_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_9_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln248_fu_1359_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TDATA_blk_n = weight_V_V_TVALID;
    end else begin
        weight_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_1359_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TREADY = 1'b1;
    end else begin
        weight_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln248_fu_1359_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((ap_enable_reg_pp0_iter3 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter3 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln248_fu_1359_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accu_0_0_V_fu_2837_p2 = ($signed(add_ln700_2_fu_2815_p2) + $signed(sext_ln700_6_fu_2833_p1));

assign accu_0_1_V_fu_2877_p2 = ($signed(add_ln700_10_fu_2855_p2) + $signed(sext_ln700_13_fu_2873_p1));

assign accu_0_2_V_fu_2917_p2 = ($signed(add_ln700_18_fu_2895_p2) + $signed(sext_ln700_20_fu_2913_p1));

assign accu_0_3_V_fu_2957_p2 = ($signed(add_ln700_26_fu_2935_p2) + $signed(sext_ln700_27_fu_2953_p1));

assign add_ln700_10_fu_2855_p2 = ($signed(add_ln700_8_fu_2846_p2) + $signed(sext_ln700_9_fu_2852_p1));

assign add_ln700_11_fu_2397_p2 = ($signed(sext_ln170_6_fu_2300_p1) + $signed(sext_ln170_9_fu_2339_p1));

assign add_ln700_12_fu_2403_p2 = ($signed(sext_ln700_8_fu_2387_p1) + $signed(sext_ln170_7_fu_2313_p1));

assign add_ln700_13_fu_2413_p2 = ($signed(sext_ln170_8_fu_2326_p1) + $signed(sext_ln700_11_fu_2409_p1));

assign add_ln700_14_fu_2867_p2 = ($signed(sext_ln700_10_fu_2861_p1) + $signed(sext_ln700_12_fu_2864_p1));

assign add_ln700_16_fu_2886_p2 = ($signed(sext_ln700_14_fu_2883_p1) + $signed(select_ln271_1_fu_2782_p3));

assign add_ln700_17_fu_2519_p2 = ($signed(sext_ln170_16_fu_2480_p1) + $signed(sext_ln170_17_fu_2502_p1));

assign add_ln700_18_fu_2895_p2 = ($signed(add_ln700_16_fu_2886_p2) + $signed(sext_ln700_16_fu_2892_p1));

assign add_ln700_19_fu_2525_p2 = ($signed(sext_ln170_12_fu_2428_p1) + $signed(sext_ln170_15_fu_2467_p1));

assign add_ln700_1_fu_2263_p2 = ($signed(sext_ln170_4_fu_2182_p1) + $signed(sext_ln170_5_fu_2232_p1));

assign add_ln700_20_fu_2531_p2 = ($signed(sext_ln700_15_fu_2515_p1) + $signed(sext_ln170_13_fu_2441_p1));

assign add_ln700_21_fu_2541_p2 = ($signed(sext_ln170_14_fu_2454_p1) + $signed(sext_ln700_18_fu_2537_p1));

assign add_ln700_22_fu_2907_p2 = ($signed(sext_ln700_17_fu_2901_p1) + $signed(sext_ln700_19_fu_2904_p1));

assign add_ln700_24_fu_2926_p2 = ($signed(sext_ln700_21_fu_2923_p1) + $signed(select_ln271_fu_2775_p3));

assign add_ln700_25_fu_2647_p2 = ($signed(sext_ln170_22_fu_2608_p1) + $signed(sext_ln170_23_fu_2630_p1));

assign add_ln700_26_fu_2935_p2 = ($signed(add_ln700_24_fu_2926_p2) + $signed(sext_ln700_23_fu_2932_p1));

assign add_ln700_27_fu_2653_p2 = ($signed(sext_ln170_18_fu_2556_p1) + $signed(sext_ln170_21_fu_2595_p1));

assign add_ln700_28_fu_2659_p2 = ($signed(sext_ln700_22_fu_2643_p1) + $signed(sext_ln170_19_fu_2569_p1));

assign add_ln700_29_fu_2669_p2 = ($signed(sext_ln170_20_fu_2582_p1) + $signed(sext_ln700_25_fu_2665_p1));

assign add_ln700_2_fu_2815_p2 = ($signed(add_ln700_fu_2806_p2) + $signed(sext_ln700_2_fu_2812_p1));

assign add_ln700_30_fu_2947_p2 = ($signed(sext_ln700_24_fu_2941_p1) + $signed(sext_ln700_26_fu_2944_p1));

assign add_ln700_32_fu_4090_p2 = (zext_ln142_1_fu_4077_p1 + zext_ln142_2_fu_4086_p1);

assign add_ln700_33_fu_4100_p2 = (zext_ln700_1_fu_4096_p1 + select_ln700_fu_4064_p3);

assign add_ln700_34_fu_3466_p2 = (zext_ln142_3_fu_3372_p1 + zext_ln142_4_fu_3381_p1);

assign add_ln700_35_fu_3476_p2 = (zext_ln142_5_fu_3390_p1 + zext_ln142_6_fu_3399_p1);

assign add_ln700_36_fu_3486_p2 = (zext_ln700_3_fu_3482_p1 + zext_ln700_2_fu_3472_p1);

assign add_ln700_37_fu_4109_p2 = (zext_ln700_4_fu_4106_p1 + add_ln700_33_fu_4100_p2);

assign add_ln700_38_fu_3492_p2 = (zext_ln142_8_fu_3417_p1 + zext_ln142_9_fu_3426_p1);

assign add_ln700_39_fu_3498_p2 = (add_ln700_38_fu_3492_p2 + zext_ln142_7_fu_3408_p1);

assign add_ln700_3_fu_2269_p2 = ($signed(sext_ln170_fu_2074_p1) + $signed(sext_ln170_3_fu_2155_p1));

assign add_ln700_40_fu_3508_p2 = (zext_ln142_10_fu_3435_p1 + zext_ln142_11_fu_3444_p1);

assign add_ln700_41_fu_3518_p2 = (zext_ln142_12_fu_3453_p1 + zext_ln700_fu_3462_p1);

assign add_ln700_42_fu_3528_p2 = (zext_ln700_7_fu_3524_p1 + zext_ln700_6_fu_3514_p1);

assign add_ln700_43_fu_3534_p2 = (add_ln700_42_fu_3528_p2 + zext_ln700_5_fu_3504_p1);

assign add_ln700_44_fu_4118_p2 = (zext_ln700_8_fu_4115_p1 + add_ln700_37_fu_4109_p2);

assign add_ln700_45_fu_4155_p2 = (zext_ln142_13_fu_4142_p1 + zext_ln142_14_fu_4151_p1);

assign add_ln700_46_fu_4165_p2 = (zext_ln700_10_fu_4161_p1 + select_ln700_1_fu_4129_p3);

assign add_ln700_47_fu_3639_p2 = (zext_ln142_15_fu_3545_p1 + zext_ln142_16_fu_3554_p1);

assign add_ln700_48_fu_3649_p2 = (zext_ln142_17_fu_3563_p1 + zext_ln142_18_fu_3572_p1);

assign add_ln700_49_fu_3659_p2 = (zext_ln700_12_fu_3655_p1 + zext_ln700_11_fu_3645_p1);

assign add_ln700_4_fu_2275_p2 = ($signed(sext_ln700_1_fu_2259_p1) + $signed(sext_ln170_1_fu_2101_p1));

assign add_ln700_50_fu_4174_p2 = (zext_ln700_13_fu_4171_p1 + add_ln700_46_fu_4165_p2);

assign add_ln700_51_fu_3665_p2 = (zext_ln142_20_fu_3590_p1 + zext_ln142_21_fu_3599_p1);

assign add_ln700_52_fu_3671_p2 = (add_ln700_51_fu_3665_p2 + zext_ln142_19_fu_3581_p1);

assign add_ln700_53_fu_3681_p2 = (zext_ln142_22_fu_3608_p1 + zext_ln142_23_fu_3617_p1);

assign add_ln700_54_fu_3691_p2 = (zext_ln142_24_fu_3626_p1 + zext_ln700_9_fu_3635_p1);

assign add_ln700_55_fu_3701_p2 = (zext_ln700_16_fu_3697_p1 + zext_ln700_15_fu_3687_p1);

assign add_ln700_56_fu_3707_p2 = (add_ln700_55_fu_3701_p2 + zext_ln700_14_fu_3677_p1);

assign add_ln700_57_fu_4183_p2 = (zext_ln700_17_fu_4180_p1 + add_ln700_50_fu_4174_p2);

assign add_ln700_58_fu_4220_p2 = (zext_ln142_25_fu_4207_p1 + zext_ln142_26_fu_4216_p1);

assign add_ln700_59_fu_4230_p2 = (zext_ln700_19_fu_4226_p1 + select_ln700_2_fu_4194_p3);

assign add_ln700_5_fu_2285_p2 = ($signed(sext_ln170_2_fu_2128_p1) + $signed(sext_ln700_4_fu_2281_p1));

assign add_ln700_60_fu_3812_p2 = (zext_ln142_27_fu_3718_p1 + zext_ln142_28_fu_3727_p1);

assign add_ln700_61_fu_3822_p2 = (zext_ln142_29_fu_3736_p1 + zext_ln142_30_fu_3745_p1);

assign add_ln700_62_fu_3832_p2 = (zext_ln700_21_fu_3828_p1 + zext_ln700_20_fu_3818_p1);

assign add_ln700_63_fu_4239_p2 = (zext_ln700_22_fu_4236_p1 + add_ln700_59_fu_4230_p2);

assign add_ln700_64_fu_3838_p2 = (zext_ln142_32_fu_3763_p1 + zext_ln142_33_fu_3772_p1);

assign add_ln700_65_fu_3844_p2 = (add_ln700_64_fu_3838_p2 + zext_ln142_31_fu_3754_p1);

assign add_ln700_66_fu_3854_p2 = (zext_ln142_34_fu_3781_p1 + zext_ln142_35_fu_3790_p1);

assign add_ln700_67_fu_3864_p2 = (zext_ln142_36_fu_3799_p1 + zext_ln700_18_fu_3808_p1);

assign add_ln700_68_fu_3874_p2 = (zext_ln700_25_fu_3870_p1 + zext_ln700_24_fu_3860_p1);

assign add_ln700_69_fu_3880_p2 = (add_ln700_68_fu_3874_p2 + zext_ln700_23_fu_3850_p1);

assign add_ln700_6_fu_2827_p2 = ($signed(sext_ln700_3_fu_2821_p1) + $signed(sext_ln700_5_fu_2824_p1));

assign add_ln700_70_fu_4248_p2 = (zext_ln700_26_fu_4245_p1 + add_ln700_63_fu_4239_p2);

assign add_ln700_71_fu_4285_p2 = (zext_ln142_37_fu_4272_p1 + zext_ln142_38_fu_4281_p1);

assign add_ln700_72_fu_4295_p2 = (zext_ln700_28_fu_4291_p1 + select_ln700_3_fu_4259_p3);

assign add_ln700_73_fu_3985_p2 = (zext_ln142_39_fu_3891_p1 + zext_ln142_40_fu_3900_p1);

assign add_ln700_74_fu_3995_p2 = (zext_ln142_41_fu_3909_p1 + zext_ln142_42_fu_3918_p1);

assign add_ln700_75_fu_4005_p2 = (zext_ln700_30_fu_4001_p1 + zext_ln700_29_fu_3991_p1);

assign add_ln700_76_fu_4304_p2 = (zext_ln700_31_fu_4301_p1 + add_ln700_72_fu_4295_p2);

assign add_ln700_77_fu_4011_p2 = (zext_ln142_44_fu_3936_p1 + zext_ln142_45_fu_3945_p1);

assign add_ln700_78_fu_4017_p2 = (add_ln700_77_fu_4011_p2 + zext_ln142_43_fu_3927_p1);

assign add_ln700_79_fu_4027_p2 = (zext_ln142_46_fu_3954_p1 + zext_ln142_47_fu_3963_p1);

assign add_ln700_80_fu_4037_p2 = (zext_ln142_48_fu_3972_p1 + zext_ln700_27_fu_3981_p1);

assign add_ln700_81_fu_4047_p2 = (zext_ln700_34_fu_4043_p1 + zext_ln700_33_fu_4033_p1);

assign add_ln700_82_fu_4053_p2 = (add_ln700_81_fu_4047_p2 + zext_ln700_32_fu_4023_p1);

assign add_ln700_83_fu_4313_p2 = (zext_ln700_35_fu_4310_p1 + add_ln700_76_fu_4304_p2);

assign add_ln700_8_fu_2846_p2 = ($signed(sext_ln700_7_fu_2843_p1) + $signed(select_ln271_2_fu_2789_p3));

assign add_ln700_9_fu_2391_p2 = ($signed(sext_ln170_10_fu_2352_p1) + $signed(sext_ln170_11_fu_2374_p1));

assign add_ln700_fu_2806_p2 = ($signed(sext_ln700_fu_2803_p1) + $signed(select_ln271_3_fu_2796_p3));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op98_read_state2 == 1'b1)) | ((icmp_ln248_fu_1359_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_block_state6_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op98_read_state2 == 1'b1)) | ((icmp_ln248_fu_1359_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_block_state6_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op98_read_state2 == 1'b1)) | ((icmp_ln248_fu_1359_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op98_read_state2 == 1'b1)) | ((icmp_ln248_fu_1359_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state6_io = ((icmp_ln289_reg_4790_pp0_iter3_reg == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_reg_pp0_iter0_act_m_val_V_reg_1278 = 'bx;

always @ (*) begin
    ap_predicate_op98_read_state2 = ((icmp_ln252_fu_1374_p2 == 1'd1) & (icmp_ln248_fu_1359_p2 == 1'd0));
end

assign arg_V_read_assign_1_fu_2078_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278[7:4]}};

assign arg_V_read_assign_2_fu_2105_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278[11:8]}};

assign arg_V_read_assign_3_fu_2132_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278[15:12]}};

assign arg_V_read_assign_4_fu_2159_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278[19:16]}};

assign arg_V_read_assign_5_fu_2186_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278[23:20]}};

assign arg_V_read_assign_6_fu_2209_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278[27:24]}};

assign arg_V_read_assign_7_fu_2236_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278[31:28]}};

assign i_fu_1365_p2 = (i_0_reg_1267 + 13'd1);

assign icmp_ln248_fu_1359_p2 = ((i_0_reg_1267 == 13'd4096) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_1374_p2 = ((ap_sig_allocacmp_nf_assign_load_1 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln271_fu_1720_p2 = ((sf_1_fu_384 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln289_fu_2046_p2 = ((sf_fu_2040_p2 == 32'd32) ? 1'b1 : 1'b0);

assign icmp_ln301_fu_2744_p2 = ((nf_fu_2738_p2 == 32'd128) ? 1'b1 : 1'b0);

assign icmp_ln899_10_fu_3051_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_53_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_11_fu_3057_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_52_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_12_fu_3063_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_51_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_13_fu_3069_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_50_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_14_fu_3075_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(threshs_m_thresholds_41_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_15_fu_3081_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(threshs_m_thresholds_40_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_16_fu_3087_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(threshs_m_thresholds_35_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_17_fu_3093_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(threshs_m_thresholds_34_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_18_fu_3103_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(sext_ln142_2_fu_3099_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_19_fu_3113_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(sext_ln142_3_fu_3109_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_1_fu_2997_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(sext_ln142_1_fu_2993_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_20_fu_3123_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(sext_ln142_4_fu_3119_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_21_fu_3133_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(sext_ln142_5_fu_3129_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_22_fu_3143_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(sext_ln142_6_fu_3139_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_23_fu_3153_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(sext_ln142_7_fu_3149_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_24_fu_3163_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(sext_ln142_8_fu_3159_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_25_fu_3173_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(sext_ln142_9_fu_3169_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_26_fu_3183_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(sext_ln142_10_fu_3179_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_27_fu_3193_p2 = (($signed(accu_0_1_V_fu_2877_p2) < $signed(sext_ln142_11_fu_3189_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_28_fu_3199_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_27_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_29_fu_3205_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_26_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_2_fu_3003_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_49_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_30_fu_3211_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_21_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_31_fu_3217_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_20_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_32_fu_3223_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_19_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_33_fu_3229_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_18_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_34_fu_3235_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_17_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_35_fu_3241_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_16_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_36_fu_3247_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_15_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_37_fu_3253_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_14_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_38_fu_3259_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_25_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_39_fu_3265_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_24_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_3_fu_3009_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_48_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_40_fu_3271_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_23_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_41_fu_3277_p2 = (($signed(accu_0_2_V_fu_2917_p2) < $signed(threshs_m_thresholds_22_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_42_fu_3283_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_13_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_43_fu_3289_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_12_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_44_fu_3295_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_7_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_45_fu_3301_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_6_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_46_fu_3307_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_5_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_47_fu_3313_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_4_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_48_fu_3319_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_3_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_49_fu_3325_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_2_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_4_fu_3015_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_47_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_50_fu_3331_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_1_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_51_fu_3337_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_52_fu_3343_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_11_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_53_fu_3349_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_10_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_54_fu_3355_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_9_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_55_fu_3361_p2 = (($signed(accu_0_3_V_fu_2957_p2) < $signed(threshs_m_thresholds_8_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_5_fu_3021_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_46_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_6_fu_3027_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_45_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_7_fu_3033_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_44_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_8_fu_3039_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_43_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_9_fu_3045_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(threshs_m_thresholds_42_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_fu_2987_p2 = (($signed(accu_0_0_V_fu_2837_p2) < $signed(sext_ln142_fu_2983_p1)) ? 1'b1 : 1'b0);

assign inElem_V_1_fu_1483_p33 = sf_1_fu_384[4:0];

assign mul_ln1352_10_fu_2320_p0 = zext_ln215_2_fu_2118_p1;

assign mul_ln1352_11_fu_2333_p0 = zext_ln215_3_fu_2145_p1;

assign mul_ln1352_12_fu_2346_p0 = zext_ln215_4_fu_2172_p1;

assign mul_ln1352_13_fu_2359_p0 = zext_ln215_5_fu_2199_p1;

assign mul_ln1352_14_fu_2368_p0 = zext_ln215_6_fu_2222_p1;

assign mul_ln1352_15_fu_2381_p0 = zext_ln215_7_fu_2249_p1;

assign mul_ln1352_16_fu_2422_p0 = zext_ln215_fu_2064_p1;

assign mul_ln1352_17_fu_2435_p0 = zext_ln215_1_fu_2091_p1;

assign mul_ln1352_18_fu_2448_p0 = zext_ln215_2_fu_2118_p1;

assign mul_ln1352_19_fu_2461_p0 = zext_ln215_3_fu_2145_p1;

assign mul_ln1352_1_fu_2095_p0 = zext_ln215_1_fu_2091_p1;

assign mul_ln1352_20_fu_2474_p0 = zext_ln215_4_fu_2172_p1;

assign mul_ln1352_21_fu_2487_p0 = zext_ln215_5_fu_2199_p1;

assign mul_ln1352_22_fu_2496_p0 = zext_ln215_6_fu_2222_p1;

assign mul_ln1352_23_fu_2509_p0 = zext_ln215_7_fu_2249_p1;

assign mul_ln1352_24_fu_2550_p0 = zext_ln215_fu_2064_p1;

assign mul_ln1352_25_fu_2563_p0 = zext_ln215_1_fu_2091_p1;

assign mul_ln1352_26_fu_2576_p0 = zext_ln215_2_fu_2118_p1;

assign mul_ln1352_27_fu_2589_p0 = zext_ln215_3_fu_2145_p1;

assign mul_ln1352_28_fu_2602_p0 = zext_ln215_4_fu_2172_p1;

assign mul_ln1352_29_fu_2615_p0 = zext_ln215_5_fu_2199_p1;

assign mul_ln1352_2_fu_2122_p0 = zext_ln215_2_fu_2118_p1;

assign mul_ln1352_30_fu_2624_p0 = zext_ln215_6_fu_2222_p1;

assign mul_ln1352_31_fu_2637_p0 = zext_ln215_7_fu_2249_p1;

assign mul_ln1352_3_fu_2149_p0 = zext_ln215_3_fu_2145_p1;

assign mul_ln1352_4_fu_2176_p0 = zext_ln215_4_fu_2172_p1;

assign mul_ln1352_5_fu_2203_p0 = zext_ln215_5_fu_2199_p1;

assign mul_ln1352_6_fu_2226_p0 = zext_ln215_6_fu_2222_p1;

assign mul_ln1352_7_fu_2253_p0 = zext_ln215_7_fu_2249_p1;

assign mul_ln1352_8_fu_2294_p0 = zext_ln215_fu_2064_p1;

assign mul_ln1352_9_fu_2307_p0 = zext_ln215_1_fu_2091_p1;

assign mul_ln1352_fu_2068_p0 = zext_ln215_fu_2064_p1;

assign nf_fu_2738_p2 = (nf_assign_fu_516 + 32'd1);

assign out_V_V_TDATA = {{{{add_ln700_83_fu_4313_p2}, {add_ln700_70_fu_4248_p2}}, {add_ln700_57_fu_4183_p2}}, {add_ln700_44_fu_4118_p2}};

assign select_ln271_1_fu_2782_p3 = ((icmp_ln271_reg_4622_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_2_0_fu_376);

assign select_ln271_2_fu_2789_p3 = ((icmp_ln271_reg_4622_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_1_0_fu_372);

assign select_ln271_3_fu_2796_p3 = ((icmp_ln271_reg_4622_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_0_0_fu_368);

assign select_ln271_fu_2775_p3 = ((icmp_ln271_reg_4622_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_3_0_fu_380);

assign select_ln301_fu_2750_p3 = ((icmp_ln301_fu_2744_p2[0:0] === 1'b1) ? 32'd0 : nf_fu_2738_p2);

assign select_ln700_1_fu_4129_p3 = ((xor_ln899_14_fu_4124_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign select_ln700_2_fu_4194_p3 = ((xor_ln899_28_fu_4189_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign select_ln700_3_fu_4259_p3 = ((xor_ln899_42_fu_4254_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign select_ln700_fu_4064_p3 = ((xor_ln899_fu_4059_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign sext_ln142_10_fu_3179_p1 = $signed(threshs_m_thresholds_37_q0);

assign sext_ln142_11_fu_3189_p1 = $signed(threshs_m_thresholds_36_q0);

assign sext_ln142_1_fu_2993_p1 = $signed(threshs_m_thresholds_54_q0);

assign sext_ln142_2_fu_3099_p1 = $signed(threshs_m_thresholds_33_q0);

assign sext_ln142_3_fu_3109_p1 = $signed(threshs_m_thresholds_32_q0);

assign sext_ln142_4_fu_3119_p1 = $signed(threshs_m_thresholds_31_q0);

assign sext_ln142_5_fu_3129_p1 = $signed(threshs_m_thresholds_30_q0);

assign sext_ln142_6_fu_3139_p1 = $signed(threshs_m_thresholds_29_q0);

assign sext_ln142_7_fu_3149_p1 = $signed(threshs_m_thresholds_28_q0);

assign sext_ln142_8_fu_3159_p1 = $signed(threshs_m_thresholds_39_q0);

assign sext_ln142_9_fu_3169_p1 = $signed(threshs_m_thresholds_38_q0);

assign sext_ln142_fu_2983_p1 = $signed(threshs_m_thresholds_55_q0);

assign sext_ln170_10_fu_2352_p1 = mul_ln1352_12_fu_2346_p2;

assign sext_ln170_11_fu_2374_p1 = mul_ln1352_14_fu_2368_p2;

assign sext_ln170_12_fu_2428_p1 = mul_ln1352_16_fu_2422_p2;

assign sext_ln170_13_fu_2441_p1 = mul_ln1352_17_fu_2435_p2;

assign sext_ln170_14_fu_2454_p1 = mul_ln1352_18_fu_2448_p2;

assign sext_ln170_15_fu_2467_p1 = mul_ln1352_19_fu_2461_p2;

assign sext_ln170_16_fu_2480_p1 = mul_ln1352_20_fu_2474_p2;

assign sext_ln170_17_fu_2502_p1 = mul_ln1352_22_fu_2496_p2;

assign sext_ln170_18_fu_2556_p1 = mul_ln1352_24_fu_2550_p2;

assign sext_ln170_19_fu_2569_p1 = mul_ln1352_25_fu_2563_p2;

assign sext_ln170_1_fu_2101_p1 = mul_ln1352_1_fu_2095_p2;

assign sext_ln170_20_fu_2582_p1 = mul_ln1352_26_fu_2576_p2;

assign sext_ln170_21_fu_2595_p1 = mul_ln1352_27_fu_2589_p2;

assign sext_ln170_22_fu_2608_p1 = mul_ln1352_28_fu_2602_p2;

assign sext_ln170_23_fu_2630_p1 = mul_ln1352_30_fu_2624_p2;

assign sext_ln170_2_fu_2128_p1 = mul_ln1352_2_fu_2122_p2;

assign sext_ln170_3_fu_2155_p1 = mul_ln1352_3_fu_2149_p2;

assign sext_ln170_4_fu_2182_p1 = mul_ln1352_4_fu_2176_p2;

assign sext_ln170_5_fu_2232_p1 = mul_ln1352_6_fu_2226_p2;

assign sext_ln170_6_fu_2300_p1 = mul_ln1352_8_fu_2294_p2;

assign sext_ln170_7_fu_2313_p1 = mul_ln1352_9_fu_2307_p2;

assign sext_ln170_8_fu_2326_p1 = mul_ln1352_10_fu_2320_p2;

assign sext_ln170_9_fu_2339_p1 = mul_ln1352_11_fu_2333_p2;

assign sext_ln170_fu_2074_p1 = mul_ln1352_fu_2068_p2;

assign sext_ln700_10_fu_2861_p1 = $signed(add_ln700_11_reg_4824);

assign sext_ln700_11_fu_2409_p1 = $signed(add_ln700_12_fu_2403_p2);

assign sext_ln700_12_fu_2864_p1 = $signed(add_ln700_13_reg_4829);

assign sext_ln700_13_fu_2873_p1 = $signed(add_ln700_14_fu_2867_p2);

assign sext_ln700_14_fu_2883_p1 = mul_ln1352_21_reg_4834;

assign sext_ln700_15_fu_2515_p1 = mul_ln1352_23_fu_2509_p2;

assign sext_ln700_16_fu_2892_p1 = $signed(add_ln700_17_reg_4839);

assign sext_ln700_17_fu_2901_p1 = $signed(add_ln700_19_reg_4844);

assign sext_ln700_18_fu_2537_p1 = $signed(add_ln700_20_fu_2531_p2);

assign sext_ln700_19_fu_2904_p1 = $signed(add_ln700_21_reg_4849);

assign sext_ln700_1_fu_2259_p1 = mul_ln1352_7_fu_2253_p2;

assign sext_ln700_20_fu_2913_p1 = $signed(add_ln700_22_fu_2907_p2);

assign sext_ln700_21_fu_2923_p1 = mul_ln1352_29_reg_4854;

assign sext_ln700_22_fu_2643_p1 = mul_ln1352_31_fu_2637_p2;

assign sext_ln700_23_fu_2932_p1 = $signed(add_ln700_25_reg_4859);

assign sext_ln700_24_fu_2941_p1 = $signed(add_ln700_27_reg_4864);

assign sext_ln700_25_fu_2665_p1 = $signed(add_ln700_28_fu_2659_p2);

assign sext_ln700_26_fu_2944_p1 = $signed(add_ln700_29_reg_4869);

assign sext_ln700_27_fu_2953_p1 = $signed(add_ln700_30_fu_2947_p2);

assign sext_ln700_2_fu_2812_p1 = $signed(add_ln700_1_reg_4799);

assign sext_ln700_3_fu_2821_p1 = $signed(add_ln700_3_reg_4804);

assign sext_ln700_4_fu_2281_p1 = $signed(add_ln700_4_fu_2275_p2);

assign sext_ln700_5_fu_2824_p1 = $signed(add_ln700_5_reg_4809);

assign sext_ln700_6_fu_2833_p1 = $signed(add_ln700_6_fu_2827_p2);

assign sext_ln700_7_fu_2843_p1 = mul_ln1352_13_reg_4814;

assign sext_ln700_8_fu_2387_p1 = mul_ln1352_15_fu_2381_p2;

assign sext_ln700_9_fu_2852_p1 = $signed(add_ln700_9_reg_4819);

assign sext_ln700_fu_2803_p1 = mul_ln1352_5_reg_4794;

assign sf_fu_2040_p2 = (32'd1 + sf_1_fu_384);

assign threshs_m_thresholds_10_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_11_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_12_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_13_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_14_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_15_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_16_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_17_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_18_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_19_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_1_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_20_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_21_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_22_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_23_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_24_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_25_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_26_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_27_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_28_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_29_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_2_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_30_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_31_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_32_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_33_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_34_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_35_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_36_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_37_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_38_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_39_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_3_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_40_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_41_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_42_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_43_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_44_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_45_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_46_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_47_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_48_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_49_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_4_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_50_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_51_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_52_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_53_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_54_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_55_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_5_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_6_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_7_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_8_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_9_address0 = zext_ln142_fu_2678_p1;

assign threshs_m_thresholds_address0 = zext_ln142_fu_2678_p1;

assign trunc_ln321_fu_1553_p1 = sf_1_fu_384[4:0];

assign trunc_ln647_fu_2057_p1 = ap_phi_reg_pp0_iter1_act_m_val_V_reg_1278[3:0];

assign wgt_M_instance_0_V_fu_1726_p1 = weight_V_V_TDATA[3:0];

assign xor_ln899_10_fu_3430_p2 = (icmp_ln899_10_reg_5204 ^ 1'd1);

assign xor_ln899_11_fu_3439_p2 = (icmp_ln899_11_reg_5209 ^ 1'd1);

assign xor_ln899_12_fu_3448_p2 = (icmp_ln899_12_reg_5214 ^ 1'd1);

assign xor_ln899_13_fu_3457_p2 = (icmp_ln899_13_reg_5219 ^ 1'd1);

assign xor_ln899_14_fu_4124_p2 = (icmp_ln899_14_reg_5224_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_15_fu_4137_p2 = (icmp_ln899_15_reg_5229_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_16_fu_4146_p2 = (icmp_ln899_16_reg_5234_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_17_fu_3540_p2 = (icmp_ln899_17_reg_5239 ^ 1'd1);

assign xor_ln899_18_fu_3549_p2 = (icmp_ln899_18_reg_5244 ^ 1'd1);

assign xor_ln899_19_fu_3558_p2 = (icmp_ln899_19_reg_5249 ^ 1'd1);

assign xor_ln899_1_fu_4072_p2 = (icmp_ln899_1_reg_5159_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_20_fu_3567_p2 = (icmp_ln899_20_reg_5254 ^ 1'd1);

assign xor_ln899_21_fu_3576_p2 = (icmp_ln899_21_reg_5259 ^ 1'd1);

assign xor_ln899_22_fu_3585_p2 = (icmp_ln899_22_reg_5264 ^ 1'd1);

assign xor_ln899_23_fu_3594_p2 = (icmp_ln899_23_reg_5269 ^ 1'd1);

assign xor_ln899_24_fu_3603_p2 = (icmp_ln899_24_reg_5274 ^ 1'd1);

assign xor_ln899_25_fu_3612_p2 = (icmp_ln899_25_reg_5279 ^ 1'd1);

assign xor_ln899_26_fu_3621_p2 = (icmp_ln899_26_reg_5284 ^ 1'd1);

assign xor_ln899_27_fu_3630_p2 = (icmp_ln899_27_reg_5289 ^ 1'd1);

assign xor_ln899_28_fu_4189_p2 = (icmp_ln899_28_reg_5294_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_29_fu_4202_p2 = (icmp_ln899_29_reg_5299_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_2_fu_4081_p2 = (icmp_ln899_2_reg_5164_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_30_fu_4211_p2 = (icmp_ln899_30_reg_5304_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_31_fu_3713_p2 = (icmp_ln899_31_reg_5309 ^ 1'd1);

assign xor_ln899_32_fu_3722_p2 = (icmp_ln899_32_reg_5314 ^ 1'd1);

assign xor_ln899_33_fu_3731_p2 = (icmp_ln899_33_reg_5319 ^ 1'd1);

assign xor_ln899_34_fu_3740_p2 = (icmp_ln899_34_reg_5324 ^ 1'd1);

assign xor_ln899_35_fu_3749_p2 = (icmp_ln899_35_reg_5329 ^ 1'd1);

assign xor_ln899_36_fu_3758_p2 = (icmp_ln899_36_reg_5334 ^ 1'd1);

assign xor_ln899_37_fu_3767_p2 = (icmp_ln899_37_reg_5339 ^ 1'd1);

assign xor_ln899_38_fu_3776_p2 = (icmp_ln899_38_reg_5344 ^ 1'd1);

assign xor_ln899_39_fu_3785_p2 = (icmp_ln899_39_reg_5349 ^ 1'd1);

assign xor_ln899_3_fu_3367_p2 = (icmp_ln899_3_reg_5169 ^ 1'd1);

assign xor_ln899_40_fu_3794_p2 = (icmp_ln899_40_reg_5354 ^ 1'd1);

assign xor_ln899_41_fu_3803_p2 = (icmp_ln899_41_reg_5359 ^ 1'd1);

assign xor_ln899_42_fu_4254_p2 = (icmp_ln899_42_reg_5364_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_43_fu_4267_p2 = (icmp_ln899_43_reg_5369_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_44_fu_4276_p2 = (icmp_ln899_44_reg_5374_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_45_fu_3886_p2 = (icmp_ln899_45_reg_5379 ^ 1'd1);

assign xor_ln899_46_fu_3895_p2 = (icmp_ln899_46_reg_5384 ^ 1'd1);

assign xor_ln899_47_fu_3904_p2 = (icmp_ln899_47_reg_5389 ^ 1'd1);

assign xor_ln899_48_fu_3913_p2 = (icmp_ln899_48_reg_5394 ^ 1'd1);

assign xor_ln899_49_fu_3922_p2 = (icmp_ln899_49_reg_5399 ^ 1'd1);

assign xor_ln899_4_fu_3376_p2 = (icmp_ln899_4_reg_5174 ^ 1'd1);

assign xor_ln899_50_fu_3931_p2 = (icmp_ln899_50_reg_5404 ^ 1'd1);

assign xor_ln899_51_fu_3940_p2 = (icmp_ln899_51_reg_5409 ^ 1'd1);

assign xor_ln899_52_fu_3949_p2 = (icmp_ln899_52_reg_5414 ^ 1'd1);

assign xor_ln899_53_fu_3958_p2 = (icmp_ln899_53_reg_5419 ^ 1'd1);

assign xor_ln899_54_fu_3967_p2 = (icmp_ln899_54_reg_5424 ^ 1'd1);

assign xor_ln899_55_fu_3976_p2 = (icmp_ln899_55_reg_5429 ^ 1'd1);

assign xor_ln899_5_fu_3385_p2 = (icmp_ln899_5_reg_5179 ^ 1'd1);

assign xor_ln899_6_fu_3394_p2 = (icmp_ln899_6_reg_5184 ^ 1'd1);

assign xor_ln899_7_fu_3403_p2 = (icmp_ln899_7_reg_5189 ^ 1'd1);

assign xor_ln899_8_fu_3412_p2 = (icmp_ln899_8_reg_5194 ^ 1'd1);

assign xor_ln899_9_fu_3421_p2 = (icmp_ln899_9_reg_5199 ^ 1'd1);

assign xor_ln899_fu_4059_p2 = (icmp_ln899_reg_5154_pp0_iter3_reg ^ 1'd1);

assign zext_ln142_10_fu_3435_p1 = xor_ln899_10_fu_3430_p2;

assign zext_ln142_11_fu_3444_p1 = xor_ln899_11_fu_3439_p2;

assign zext_ln142_12_fu_3453_p1 = xor_ln899_12_fu_3448_p2;

assign zext_ln142_13_fu_4142_p1 = xor_ln899_15_fu_4137_p2;

assign zext_ln142_14_fu_4151_p1 = xor_ln899_16_fu_4146_p2;

assign zext_ln142_15_fu_3545_p1 = xor_ln899_17_fu_3540_p2;

assign zext_ln142_16_fu_3554_p1 = xor_ln899_18_fu_3549_p2;

assign zext_ln142_17_fu_3563_p1 = xor_ln899_19_fu_3558_p2;

assign zext_ln142_18_fu_3572_p1 = xor_ln899_20_fu_3567_p2;

assign zext_ln142_19_fu_3581_p1 = xor_ln899_21_fu_3576_p2;

assign zext_ln142_1_fu_4077_p1 = xor_ln899_1_fu_4072_p2;

assign zext_ln142_20_fu_3590_p1 = xor_ln899_22_fu_3585_p2;

assign zext_ln142_21_fu_3599_p1 = xor_ln899_23_fu_3594_p2;

assign zext_ln142_22_fu_3608_p1 = xor_ln899_24_fu_3603_p2;

assign zext_ln142_23_fu_3617_p1 = xor_ln899_25_fu_3612_p2;

assign zext_ln142_24_fu_3626_p1 = xor_ln899_26_fu_3621_p2;

assign zext_ln142_25_fu_4207_p1 = xor_ln899_29_fu_4202_p2;

assign zext_ln142_26_fu_4216_p1 = xor_ln899_30_fu_4211_p2;

assign zext_ln142_27_fu_3718_p1 = xor_ln899_31_fu_3713_p2;

assign zext_ln142_28_fu_3727_p1 = xor_ln899_32_fu_3722_p2;

assign zext_ln142_29_fu_3736_p1 = xor_ln899_33_fu_3731_p2;

assign zext_ln142_2_fu_4086_p1 = xor_ln899_2_fu_4081_p2;

assign zext_ln142_30_fu_3745_p1 = xor_ln899_34_fu_3740_p2;

assign zext_ln142_31_fu_3754_p1 = xor_ln899_35_fu_3749_p2;

assign zext_ln142_32_fu_3763_p1 = xor_ln899_36_fu_3758_p2;

assign zext_ln142_33_fu_3772_p1 = xor_ln899_37_fu_3767_p2;

assign zext_ln142_34_fu_3781_p1 = xor_ln899_38_fu_3776_p2;

assign zext_ln142_35_fu_3790_p1 = xor_ln899_39_fu_3785_p2;

assign zext_ln142_36_fu_3799_p1 = xor_ln899_40_fu_3794_p2;

assign zext_ln142_37_fu_4272_p1 = xor_ln899_43_fu_4267_p2;

assign zext_ln142_38_fu_4281_p1 = xor_ln899_44_fu_4276_p2;

assign zext_ln142_39_fu_3891_p1 = xor_ln899_45_fu_3886_p2;

assign zext_ln142_3_fu_3372_p1 = xor_ln899_3_fu_3367_p2;

assign zext_ln142_40_fu_3900_p1 = xor_ln899_46_fu_3895_p2;

assign zext_ln142_41_fu_3909_p1 = xor_ln899_47_fu_3904_p2;

assign zext_ln142_42_fu_3918_p1 = xor_ln899_48_fu_3913_p2;

assign zext_ln142_43_fu_3927_p1 = xor_ln899_49_fu_3922_p2;

assign zext_ln142_44_fu_3936_p1 = xor_ln899_50_fu_3931_p2;

assign zext_ln142_45_fu_3945_p1 = xor_ln899_51_fu_3940_p2;

assign zext_ln142_46_fu_3954_p1 = xor_ln899_52_fu_3949_p2;

assign zext_ln142_47_fu_3963_p1 = xor_ln899_53_fu_3958_p2;

assign zext_ln142_48_fu_3972_p1 = xor_ln899_54_fu_3967_p2;

assign zext_ln142_4_fu_3381_p1 = xor_ln899_4_fu_3376_p2;

assign zext_ln142_5_fu_3390_p1 = xor_ln899_5_fu_3385_p2;

assign zext_ln142_6_fu_3399_p1 = xor_ln899_6_fu_3394_p2;

assign zext_ln142_7_fu_3408_p1 = xor_ln899_7_fu_3403_p2;

assign zext_ln142_8_fu_3417_p1 = xor_ln899_8_fu_3412_p2;

assign zext_ln142_9_fu_3426_p1 = xor_ln899_9_fu_3421_p2;

assign zext_ln142_fu_2678_p1 = nf_assign_fu_516;

assign zext_ln215_1_fu_2091_p1 = arg_V_read_assign_1_fu_2078_p4;

assign zext_ln215_2_fu_2118_p1 = arg_V_read_assign_2_fu_2105_p4;

assign zext_ln215_3_fu_2145_p1 = arg_V_read_assign_3_fu_2132_p4;

assign zext_ln215_4_fu_2172_p1 = arg_V_read_assign_4_fu_2159_p4;

assign zext_ln215_5_fu_2199_p1 = arg_V_read_assign_5_fu_2186_p4;

assign zext_ln215_6_fu_2222_p1 = arg_V_read_assign_6_fu_2209_p4;

assign zext_ln215_7_fu_2249_p1 = arg_V_read_assign_7_fu_2236_p4;

assign zext_ln215_fu_2064_p1 = trunc_ln647_fu_2057_p1;

assign zext_ln700_10_fu_4161_p1 = add_ln700_45_fu_4155_p2;

assign zext_ln700_11_fu_3645_p1 = add_ln700_47_fu_3639_p2;

assign zext_ln700_12_fu_3655_p1 = add_ln700_48_fu_3649_p2;

assign zext_ln700_13_fu_4171_p1 = add_ln700_49_reg_5444;

assign zext_ln700_14_fu_3677_p1 = add_ln700_52_fu_3671_p2;

assign zext_ln700_15_fu_3687_p1 = add_ln700_53_fu_3681_p2;

assign zext_ln700_16_fu_3697_p1 = add_ln700_54_fu_3691_p2;

assign zext_ln700_17_fu_4180_p1 = add_ln700_56_reg_5449;

assign zext_ln700_18_fu_3808_p1 = xor_ln899_41_fu_3803_p2;

assign zext_ln700_19_fu_4226_p1 = add_ln700_58_fu_4220_p2;

assign zext_ln700_1_fu_4096_p1 = add_ln700_32_fu_4090_p2;

assign zext_ln700_20_fu_3818_p1 = add_ln700_60_fu_3812_p2;

assign zext_ln700_21_fu_3828_p1 = add_ln700_61_fu_3822_p2;

assign zext_ln700_22_fu_4236_p1 = add_ln700_62_reg_5454;

assign zext_ln700_23_fu_3850_p1 = add_ln700_65_fu_3844_p2;

assign zext_ln700_24_fu_3860_p1 = add_ln700_66_fu_3854_p2;

assign zext_ln700_25_fu_3870_p1 = add_ln700_67_fu_3864_p2;

assign zext_ln700_26_fu_4245_p1 = add_ln700_69_reg_5459;

assign zext_ln700_27_fu_3981_p1 = xor_ln899_55_fu_3976_p2;

assign zext_ln700_28_fu_4291_p1 = add_ln700_71_fu_4285_p2;

assign zext_ln700_29_fu_3991_p1 = add_ln700_73_fu_3985_p2;

assign zext_ln700_2_fu_3472_p1 = add_ln700_34_fu_3466_p2;

assign zext_ln700_30_fu_4001_p1 = add_ln700_74_fu_3995_p2;

assign zext_ln700_31_fu_4301_p1 = add_ln700_75_reg_5464;

assign zext_ln700_32_fu_4023_p1 = add_ln700_78_fu_4017_p2;

assign zext_ln700_33_fu_4033_p1 = add_ln700_79_fu_4027_p2;

assign zext_ln700_34_fu_4043_p1 = add_ln700_80_fu_4037_p2;

assign zext_ln700_35_fu_4310_p1 = add_ln700_82_reg_5469;

assign zext_ln700_3_fu_3482_p1 = add_ln700_35_fu_3476_p2;

assign zext_ln700_4_fu_4106_p1 = add_ln700_36_reg_5434;

assign zext_ln700_5_fu_3504_p1 = add_ln700_39_fu_3498_p2;

assign zext_ln700_6_fu_3514_p1 = add_ln700_40_fu_3508_p2;

assign zext_ln700_7_fu_3524_p1 = add_ln700_41_fu_3518_p2;

assign zext_ln700_8_fu_4115_p1 = add_ln700_43_reg_5439;

assign zext_ln700_9_fu_3635_p1 = xor_ln899_27_fu_3630_p2;

assign zext_ln700_fu_3462_p1 = xor_ln899_13_fu_3457_p2;

endmodule //StreamingFCLayer_Batch_3_Matrix_Vector_Activa
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/bc91/hdl/verilog/StreamingFCLayer_Batch_6_StreamingFCLayer_Batch_6.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingFCLayer_Batch_6_StreamingFCLayer_Batch_6,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.336000,HLS_SYN_LAT=1797,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=2167,HLS_SYN_LUT=1847,HLS_VERSION=2020_1_1}" *)

module StreamingFCLayer_Batch_6_StreamingFCLayer_Batch_6 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        weights_V_V_TDATA,
        weights_V_V_TVALID,
        weights_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [7:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
input  [7:0] weights_V_V_TDATA;
input   weights_V_V_TVALID;
output   weights_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;
reg weights_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_Matrix_Vector_Activa_fu_28_ap_start;
wire    grp_Matrix_Vector_Activa_fu_28_ap_done;
wire    grp_Matrix_Vector_Activa_fu_28_ap_idle;
wire    grp_Matrix_Vector_Activa_fu_28_ap_ready;
wire    grp_Matrix_Vector_Activa_fu_28_in_V_V_TREADY;
wire   [15:0] grp_Matrix_Vector_Activa_fu_28_out_V_V_TDATA;
wire    grp_Matrix_Vector_Activa_fu_28_out_V_V_TVALID;
wire    grp_Matrix_Vector_Activa_fu_28_out_V_V_TREADY;
wire    grp_Matrix_Vector_Activa_fu_28_weight_V_V_TREADY;
reg    grp_Matrix_Vector_Activa_fu_28_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [7:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    regslice_both_weights_V_V_U_apdone_blk;
wire   [7:0] weights_V_V_TDATA_int;
wire    weights_V_V_TVALID_int;
reg    weights_V_V_TREADY_int;
wire    regslice_both_weights_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_Matrix_Vector_Activa_fu_28_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingFCLayer_Batch_6_Matrix_Vector_Activa grp_Matrix_Vector_Activa_fu_28(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_Matrix_Vector_Activa_fu_28_ap_start),
    .ap_done(grp_Matrix_Vector_Activa_fu_28_ap_done),
    .ap_idle(grp_Matrix_Vector_Activa_fu_28_ap_idle),
    .ap_ready(grp_Matrix_Vector_Activa_fu_28_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_Matrix_Vector_Activa_fu_28_in_V_V_TREADY),
    .out_V_V_TDATA(grp_Matrix_Vector_Activa_fu_28_out_V_V_TDATA),
    .out_V_V_TVALID(grp_Matrix_Vector_Activa_fu_28_out_V_V_TVALID),
    .out_V_V_TREADY(grp_Matrix_Vector_Activa_fu_28_out_V_V_TREADY),
    .weight_V_V_TDATA(weights_V_V_TDATA_int),
    .weight_V_V_TVALID(weights_V_V_TVALID_int),
    .weight_V_V_TREADY(grp_Matrix_Vector_Activa_fu_28_weight_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_weights_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(weights_V_V_TDATA),
    .vld_in(weights_V_V_TVALID),
    .ack_in(regslice_both_weights_V_V_U_ack_in),
    .data_out(weights_V_V_TDATA_int),
    .vld_out(weights_V_V_TVALID_int),
    .ack_out(weights_V_V_TREADY_int),
    .apdone_blk(regslice_both_weights_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_Matrix_Vector_Activa_fu_28_out_V_V_TDATA),
    .vld_in(grp_Matrix_Vector_Activa_fu_28_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_Matrix_Vector_Activa_fu_28_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_Matrix_Vector_Activa_fu_28_ap_start_reg <= 1'b1;
        end else if ((grp_Matrix_Vector_Activa_fu_28_ap_ready == 1'b1)) begin
            grp_Matrix_Vector_Activa_fu_28_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_28_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    if (((regslice_both_weights_V_V_U_ack_in == 1'b1) & (weights_V_V_TVALID == 1'b1))) begin
        weights_V_V_TREADY = 1'b1;
    end else begin
        weights_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        weights_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_28_weight_V_V_TREADY;
    end else begin
        weights_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_Matrix_Vector_Activa_fu_28_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_Matrix_Vector_Activa_fu_28_ap_start = grp_Matrix_Vector_Activa_fu_28_ap_start_reg;

assign grp_Matrix_Vector_Activa_fu_28_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingFCLayer_Batch_6_StreamingFCLayer_Batch_6
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActlbW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActlbW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActlbW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActlbW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActlbW_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActlbW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActZio.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActZio_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActZio_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActZio(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActZio_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActZio_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbvn.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbvn_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbvn_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbvn(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbvn_rom Thresholding_Batch_0_Thresholding_Batcbvn_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbxn.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbxn_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbxn_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbxn(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbxn_rom Thresholding_Batch_0_Thresholding_Batcbxn_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_7_0/synth/finn_design_StreamingFIFO_7_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_7:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_7,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_7_0,StreamingFIFO_7,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_7_0,StreamingFIFO_7,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_7,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_7_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [23 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 3, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [23 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 3, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_7 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/b054/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccmv.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccmv_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccmv_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccmv(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccmv_rom Thresholding_Batch_0_Thresholding_Batccmv_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActShg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActShg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActShg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActShg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActShg_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActShg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actibs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actibs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actibs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actibs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actibs_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actibs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_1_0/synth/finn_design_StreamingFCLayer_Batch_1_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFCLayer_Batch_1:1.0
// IP Revision: 2101301320

(* X_CORE_INFO = "StreamingFCLayer_Batch_1_StreamingFCLayer_Batch_1,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_1_0,StreamingFCLayer_Batch_1_StreamingFCLayer_Batch_1,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_1_0,StreamingFCLayer_Batch_1_StreamingFCLayer_Batch_1,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFCLayer_Batch_1,x_ipVersion=1.0,x_ipCoreRevision=2101301320,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_1_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  weights_V_V_TVALID,
  weights_V_V_TREADY,
  weights_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:weights_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TVALID" *)
input wire weights_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TREADY" *)
output wire weights_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME weights_V_V, TDATA_NUM_BYTES 8, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TDATA" *)
input wire [63 : 0] weights_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;

  StreamingFCLayer_Batch_1_StreamingFCLayer_Batch_1 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .weights_V_V_TVALID(weights_V_V_TVALID),
    .weights_V_V_TREADY(weights_V_V_TREADY),
    .weights_V_V_TDATA(weights_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/e03c/hdl/verilog/ConvolutionInputGenerator_3_ConvolutionInputGbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module ConvolutionInputGenerator_3_ConvolutionInputGbkb_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 32;
parameter AWIDTH = 8;
parameter MEM_SIZE = 240;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];




always @(posedge clk)  
begin 
    if (ce0) begin
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module ConvolutionInputGenerator_3_ConvolutionInputGbkb(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd32;
parameter AddressRange = 32'd240;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



ConvolutionInputGenerator_3_ConvolutionInputGbkb_ram ConvolutionInputGenerator_3_ConvolutionInputGbkb_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActlbW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActlbW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActlbW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActlbW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActlbW_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActlbW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdcE.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcdcE_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdcE_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcdcE(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcdcE_rom Thresholding_Batch_0_Thresholding_BatcdcE_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/6405/hdl/verilog/StreamingFCLayer_Batch_5_StreamingFCLayer_bkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module StreamingFCLayer_Batch_5_StreamingFCLayer_bkb #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH       = 32,
    din5_WIDTH       = 32,
    din6_WIDTH       = 32,
    din7_WIDTH       = 32,
    din8_WIDTH       = 32,
    din9_WIDTH       = 32,
    din10_WIDTH       = 32,
    din11_WIDTH       = 32,
    din12_WIDTH       = 32,
    din13_WIDTH       = 32,
    din14_WIDTH       = 32,
    din15_WIDTH       = 32,
    din16_WIDTH       = 32,
    din17_WIDTH       = 32,
    din18_WIDTH       = 32,
    din19_WIDTH       = 32,
    din20_WIDTH       = 32,
    din21_WIDTH       = 32,
    din22_WIDTH       = 32,
    din23_WIDTH       = 32,
    din24_WIDTH       = 32,
    din25_WIDTH       = 32,
    din26_WIDTH       = 32,
    din27_WIDTH       = 32,
    din28_WIDTH       = 32,
    din29_WIDTH       = 32,
    din30_WIDTH       = 32,
    din31_WIDTH       = 32,
    din32_WIDTH       = 32,
    din33_WIDTH       = 32,
    din34_WIDTH       = 32,
    din35_WIDTH       = 32,
    din36_WIDTH       = 32,
    din37_WIDTH       = 32,
    din38_WIDTH       = 32,
    din39_WIDTH       = 32,
    din40_WIDTH       = 32,
    din41_WIDTH       = 32,
    din42_WIDTH       = 32,
    din43_WIDTH       = 32,
    din44_WIDTH       = 32,
    din45_WIDTH       = 32,
    din46_WIDTH       = 32,
    din47_WIDTH       = 32,
    din48_WIDTH       = 32,
    din49_WIDTH       = 32,
    din50_WIDTH       = 32,
    din51_WIDTH       = 32,
    din52_WIDTH       = 32,
    din53_WIDTH       = 32,
    din54_WIDTH       = 32,
    din55_WIDTH       = 32,
    din56_WIDTH       = 32,
    din57_WIDTH       = 32,
    din58_WIDTH       = 32,
    din59_WIDTH       = 32,
    din60_WIDTH       = 32,
    din61_WIDTH       = 32,
    din62_WIDTH       = 32,
    din63_WIDTH       = 32,
    din64_WIDTH       = 32,
    din65_WIDTH       = 32,
    din66_WIDTH       = 32,
    din67_WIDTH       = 32,
    din68_WIDTH       = 32,
    din69_WIDTH       = 32,
    din70_WIDTH       = 32,
    din71_WIDTH       = 32,
    din72_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [31 : 0]     din0,
    input  [31 : 0]     din1,
    input  [31 : 0]     din2,
    input  [31 : 0]     din3,
    input  [31 : 0]     din4,
    input  [31 : 0]     din5,
    input  [31 : 0]     din6,
    input  [31 : 0]     din7,
    input  [31 : 0]     din8,
    input  [31 : 0]     din9,
    input  [31 : 0]     din10,
    input  [31 : 0]     din11,
    input  [31 : 0]     din12,
    input  [31 : 0]     din13,
    input  [31 : 0]     din14,
    input  [31 : 0]     din15,
    input  [31 : 0]     din16,
    input  [31 : 0]     din17,
    input  [31 : 0]     din18,
    input  [31 : 0]     din19,
    input  [31 : 0]     din20,
    input  [31 : 0]     din21,
    input  [31 : 0]     din22,
    input  [31 : 0]     din23,
    input  [31 : 0]     din24,
    input  [31 : 0]     din25,
    input  [31 : 0]     din26,
    input  [31 : 0]     din27,
    input  [31 : 0]     din28,
    input  [31 : 0]     din29,
    input  [31 : 0]     din30,
    input  [31 : 0]     din31,
    input  [31 : 0]     din32,
    input  [31 : 0]     din33,
    input  [31 : 0]     din34,
    input  [31 : 0]     din35,
    input  [31 : 0]     din36,
    input  [31 : 0]     din37,
    input  [31 : 0]     din38,
    input  [31 : 0]     din39,
    input  [31 : 0]     din40,
    input  [31 : 0]     din41,
    input  [31 : 0]     din42,
    input  [31 : 0]     din43,
    input  [31 : 0]     din44,
    input  [31 : 0]     din45,
    input  [31 : 0]     din46,
    input  [31 : 0]     din47,
    input  [31 : 0]     din48,
    input  [31 : 0]     din49,
    input  [31 : 0]     din50,
    input  [31 : 0]     din51,
    input  [31 : 0]     din52,
    input  [31 : 0]     din53,
    input  [31 : 0]     din54,
    input  [31 : 0]     din55,
    input  [31 : 0]     din56,
    input  [31 : 0]     din57,
    input  [31 : 0]     din58,
    input  [31 : 0]     din59,
    input  [31 : 0]     din60,
    input  [31 : 0]     din61,
    input  [31 : 0]     din62,
    input  [31 : 0]     din63,
    input  [31 : 0]     din64,
    input  [31 : 0]     din65,
    input  [31 : 0]     din66,
    input  [31 : 0]     din67,
    input  [31 : 0]     din68,
    input  [31 : 0]     din69,
    input  [31 : 0]     din70,
    input  [31 : 0]     din71,
    input  [6 : 0]    din72,
    output [31 : 0]   dout);

// puts internal signals
wire [6 : 0]     sel;
// level 1 signals
wire [31 : 0]         mux_1_0;
wire [31 : 0]         mux_1_1;
wire [31 : 0]         mux_1_2;
wire [31 : 0]         mux_1_3;
wire [31 : 0]         mux_1_4;
wire [31 : 0]         mux_1_5;
wire [31 : 0]         mux_1_6;
wire [31 : 0]         mux_1_7;
wire [31 : 0]         mux_1_8;
wire [31 : 0]         mux_1_9;
wire [31 : 0]         mux_1_10;
wire [31 : 0]         mux_1_11;
wire [31 : 0]         mux_1_12;
wire [31 : 0]         mux_1_13;
wire [31 : 0]         mux_1_14;
wire [31 : 0]         mux_1_15;
wire [31 : 0]         mux_1_16;
wire [31 : 0]         mux_1_17;
wire [31 : 0]         mux_1_18;
wire [31 : 0]         mux_1_19;
wire [31 : 0]         mux_1_20;
wire [31 : 0]         mux_1_21;
wire [31 : 0]         mux_1_22;
wire [31 : 0]         mux_1_23;
wire [31 : 0]         mux_1_24;
wire [31 : 0]         mux_1_25;
wire [31 : 0]         mux_1_26;
wire [31 : 0]         mux_1_27;
wire [31 : 0]         mux_1_28;
wire [31 : 0]         mux_1_29;
wire [31 : 0]         mux_1_30;
wire [31 : 0]         mux_1_31;
wire [31 : 0]         mux_1_32;
wire [31 : 0]         mux_1_33;
wire [31 : 0]         mux_1_34;
wire [31 : 0]         mux_1_35;
// level 2 signals
wire [31 : 0]         mux_2_0;
wire [31 : 0]         mux_2_1;
wire [31 : 0]         mux_2_2;
wire [31 : 0]         mux_2_3;
wire [31 : 0]         mux_2_4;
wire [31 : 0]         mux_2_5;
wire [31 : 0]         mux_2_6;
wire [31 : 0]         mux_2_7;
wire [31 : 0]         mux_2_8;
wire [31 : 0]         mux_2_9;
wire [31 : 0]         mux_2_10;
wire [31 : 0]         mux_2_11;
wire [31 : 0]         mux_2_12;
wire [31 : 0]         mux_2_13;
wire [31 : 0]         mux_2_14;
wire [31 : 0]         mux_2_15;
wire [31 : 0]         mux_2_16;
wire [31 : 0]         mux_2_17;
// level 3 signals
wire [31 : 0]         mux_3_0;
wire [31 : 0]         mux_3_1;
wire [31 : 0]         mux_3_2;
wire [31 : 0]         mux_3_3;
wire [31 : 0]         mux_3_4;
wire [31 : 0]         mux_3_5;
wire [31 : 0]         mux_3_6;
wire [31 : 0]         mux_3_7;
wire [31 : 0]         mux_3_8;
// level 4 signals
wire [31 : 0]         mux_4_0;
wire [31 : 0]         mux_4_1;
wire [31 : 0]         mux_4_2;
wire [31 : 0]         mux_4_3;
wire [31 : 0]         mux_4_4;
// level 5 signals
wire [31 : 0]         mux_5_0;
wire [31 : 0]         mux_5_1;
wire [31 : 0]         mux_5_2;
// level 6 signals
wire [31 : 0]         mux_6_0;
wire [31 : 0]         mux_6_1;
// level 7 signals
wire [31 : 0]         mux_7_0;

assign sel = din72;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;
assign mux_1_2 = (sel[0] == 0)? din4 : din5;
assign mux_1_3 = (sel[0] == 0)? din6 : din7;
assign mux_1_4 = (sel[0] == 0)? din8 : din9;
assign mux_1_5 = (sel[0] == 0)? din10 : din11;
assign mux_1_6 = (sel[0] == 0)? din12 : din13;
assign mux_1_7 = (sel[0] == 0)? din14 : din15;
assign mux_1_8 = (sel[0] == 0)? din16 : din17;
assign mux_1_9 = (sel[0] == 0)? din18 : din19;
assign mux_1_10 = (sel[0] == 0)? din20 : din21;
assign mux_1_11 = (sel[0] == 0)? din22 : din23;
assign mux_1_12 = (sel[0] == 0)? din24 : din25;
assign mux_1_13 = (sel[0] == 0)? din26 : din27;
assign mux_1_14 = (sel[0] == 0)? din28 : din29;
assign mux_1_15 = (sel[0] == 0)? din30 : din31;
assign mux_1_16 = (sel[0] == 0)? din32 : din33;
assign mux_1_17 = (sel[0] == 0)? din34 : din35;
assign mux_1_18 = (sel[0] == 0)? din36 : din37;
assign mux_1_19 = (sel[0] == 0)? din38 : din39;
assign mux_1_20 = (sel[0] == 0)? din40 : din41;
assign mux_1_21 = (sel[0] == 0)? din42 : din43;
assign mux_1_22 = (sel[0] == 0)? din44 : din45;
assign mux_1_23 = (sel[0] == 0)? din46 : din47;
assign mux_1_24 = (sel[0] == 0)? din48 : din49;
assign mux_1_25 = (sel[0] == 0)? din50 : din51;
assign mux_1_26 = (sel[0] == 0)? din52 : din53;
assign mux_1_27 = (sel[0] == 0)? din54 : din55;
assign mux_1_28 = (sel[0] == 0)? din56 : din57;
assign mux_1_29 = (sel[0] == 0)? din58 : din59;
assign mux_1_30 = (sel[0] == 0)? din60 : din61;
assign mux_1_31 = (sel[0] == 0)? din62 : din63;
assign mux_1_32 = (sel[0] == 0)? din64 : din65;
assign mux_1_33 = (sel[0] == 0)? din66 : din67;
assign mux_1_34 = (sel[0] == 0)? din68 : din69;
assign mux_1_35 = (sel[0] == 0)? din70 : din71;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;
assign mux_2_1 = (sel[1] == 0)? mux_1_2 : mux_1_3;
assign mux_2_2 = (sel[1] == 0)? mux_1_4 : mux_1_5;
assign mux_2_3 = (sel[1] == 0)? mux_1_6 : mux_1_7;
assign mux_2_4 = (sel[1] == 0)? mux_1_8 : mux_1_9;
assign mux_2_5 = (sel[1] == 0)? mux_1_10 : mux_1_11;
assign mux_2_6 = (sel[1] == 0)? mux_1_12 : mux_1_13;
assign mux_2_7 = (sel[1] == 0)? mux_1_14 : mux_1_15;
assign mux_2_8 = (sel[1] == 0)? mux_1_16 : mux_1_17;
assign mux_2_9 = (sel[1] == 0)? mux_1_18 : mux_1_19;
assign mux_2_10 = (sel[1] == 0)? mux_1_20 : mux_1_21;
assign mux_2_11 = (sel[1] == 0)? mux_1_22 : mux_1_23;
assign mux_2_12 = (sel[1] == 0)? mux_1_24 : mux_1_25;
assign mux_2_13 = (sel[1] == 0)? mux_1_26 : mux_1_27;
assign mux_2_14 = (sel[1] == 0)? mux_1_28 : mux_1_29;
assign mux_2_15 = (sel[1] == 0)? mux_1_30 : mux_1_31;
assign mux_2_16 = (sel[1] == 0)? mux_1_32 : mux_1_33;
assign mux_2_17 = (sel[1] == 0)? mux_1_34 : mux_1_35;

// Generate level 3 logic
assign mux_3_0 = (sel[2] == 0)? mux_2_0 : mux_2_1;
assign mux_3_1 = (sel[2] == 0)? mux_2_2 : mux_2_3;
assign mux_3_2 = (sel[2] == 0)? mux_2_4 : mux_2_5;
assign mux_3_3 = (sel[2] == 0)? mux_2_6 : mux_2_7;
assign mux_3_4 = (sel[2] == 0)? mux_2_8 : mux_2_9;
assign mux_3_5 = (sel[2] == 0)? mux_2_10 : mux_2_11;
assign mux_3_6 = (sel[2] == 0)? mux_2_12 : mux_2_13;
assign mux_3_7 = (sel[2] == 0)? mux_2_14 : mux_2_15;
assign mux_3_8 = (sel[2] == 0)? mux_2_16 : mux_2_17;

// Generate level 4 logic
assign mux_4_0 = (sel[3] == 0)? mux_3_0 : mux_3_1;
assign mux_4_1 = (sel[3] == 0)? mux_3_2 : mux_3_3;
assign mux_4_2 = (sel[3] == 0)? mux_3_4 : mux_3_5;
assign mux_4_3 = (sel[3] == 0)? mux_3_6 : mux_3_7;
assign mux_4_4 = mux_3_8;

// Generate level 5 logic
assign mux_5_0 = (sel[4] == 0)? mux_4_0 : mux_4_1;
assign mux_5_1 = (sel[4] == 0)? mux_4_2 : mux_4_3;
assign mux_5_2 = mux_4_4;

// Generate level 6 logic
assign mux_6_0 = (sel[5] == 0)? mux_5_0 : mux_5_1;
assign mux_6_1 = mux_5_2;

// Generate level 7 logic
assign mux_7_0 = (sel[6] == 0)? mux_6_0 : mux_6_1;

// output logic
assign dout = mux_7_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActwdI.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActwdI_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActwdI_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActwdI(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActwdI_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActwdI_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_0_0/synth/finn_design_StreamingFCLayer_Batch_0_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFCLayer_Batch_0:1.0
// IP Revision: 2101301320

(* X_CORE_INFO = "StreamingFCLayer_Batch_0_StreamingFCLayer_Batch_0,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_0_0,StreamingFCLayer_Batch_0_StreamingFCLayer_Batch_0,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_0_0,StreamingFCLayer_Batch_0_StreamingFCLayer_Batch_0,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFCLayer_Batch_0,x_ipVersion=1.0,x_ipCoreRevision=2101301320,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_0_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  weights_V_V_TVALID,
  weights_V_V_TREADY,
  weights_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:weights_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [7 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TVALID" *)
input wire weights_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TREADY" *)
output wire weights_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME weights_V_V, TDATA_NUM_BYTES 4, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TDATA" *)
input wire [31 : 0] weights_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 12, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [95 : 0] out_V_V_TDATA;

  StreamingFCLayer_Batch_0_StreamingFCLayer_Batch_0 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .weights_V_V_TVALID(weights_V_V_TVALID),
    .weights_V_V_TREADY(weights_V_V_TREADY),
    .weights_V_V_TDATA(weights_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/2c22/hdl/verilog/ConvolutionInputGenerator_2_ConvolutionInputGenerator_2.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="ConvolutionInputGenerator_2_ConvolutionInputGenerator_2,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.027750,HLS_SYN_LAT=8201,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=540,HLS_SYN_LUT=1364,HLS_VERSION=2020_1_1}" *)

module ConvolutionInputGenerator_2_ConvolutionInputGenerator_2 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [23:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [23:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_ConvolutionInputGene_1_fu_26_ap_start;
wire    grp_ConvolutionInputGene_1_fu_26_ap_done;
wire    grp_ConvolutionInputGene_1_fu_26_ap_idle;
wire    grp_ConvolutionInputGene_1_fu_26_ap_ready;
wire    grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY;
wire   [23:0] grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA;
wire    grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID;
wire    grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY;
reg    grp_ConvolutionInputGene_1_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [23:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_ConvolutionInputGene_1_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

ConvolutionInputGenerator_2_ConvolutionInputGene_1 grp_ConvolutionInputGene_1_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_ConvolutionInputGene_1_fu_26_ap_start),
    .ap_done(grp_ConvolutionInputGene_1_fu_26_ap_done),
    .ap_idle(grp_ConvolutionInputGene_1_fu_26_ap_idle),
    .ap_ready(grp_ConvolutionInputGene_1_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 24 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 24 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA),
    .vld_in(grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_ConvolutionInputGene_1_fu_26_ap_ready == 1'b1)) begin
            grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_ConvolutionInputGene_1_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_ConvolutionInputGene_1_fu_26_ap_start = grp_ConvolutionInputGene_1_fu_26_ap_start_reg;

assign grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //ConvolutionInputGenerator_2_ConvolutionInputGenerator_2
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActJfO.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActJfO_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActJfO_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActJfO(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActJfO_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActJfO_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccsw.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccsw_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccsw_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccsw(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccsw_rom Thresholding_Batch_0_Thresholding_Batccsw_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_ConvolutionInputGenerator_1_0/synth/finn_design_ConvolutionInputGenerator_1_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:ConvolutionInputGenerator_1:1.0
// IP Revision: 2101301318

(* X_CORE_INFO = "ConvolutionInputGenerator_1_ConvolutionInputGenerator_1,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_ConvolutionInputGenerator_1_0,ConvolutionInputGenerator_1_ConvolutionInputGenerator_1,{}" *)
(* CORE_GENERATION_INFO = "finn_design_ConvolutionInputGenerator_1_0,ConvolutionInputGenerator_1_ConvolutionInputGenerator_1,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=ConvolutionInputGenerator_1,x_ipVersion=1.0,x_ipCoreRevision=2101301318,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_ConvolutionInputGenerator_1_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;

  ConvolutionInputGenerator_1_ConvolutionInputGenerator_1 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/32c2/hdl/verilog/StreamingDataWidthConverter_Batch_5_StreamingDataWidthCo_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingDataWidthConverter_Batch_5_StreamingDataWidthCo_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [15:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln370_fu_104_p2;
wire   [0:0] icmp_ln373_fu_116_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln370_reg_162;
reg   [7:0] p_025_0_reg_61;
reg   [31:0] o_0_reg_73;
reg   [8:0] t_0_reg_84;
reg    ap_predicate_op16_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [8:0] t_fu_110_p2;
reg   [0:0] icmp_ln373_reg_171;
wire   [31:0] select_ln384_fu_134_p3;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg   [15:0] ap_phi_mux_p_Val2_s_phi_fu_98_p4;
wire   [15:0] ap_phi_reg_pp0_iter0_p_Val2_s_reg_95;
reg   [15:0] ap_phi_reg_pp0_iter1_p_Val2_s_reg_95;
wire   [15:0] zext_ln370_fu_142_p1;
reg    ap_block_pp0_stage0_01001;
wire   [31:0] o_fu_122_p2;
wire   [0:0] icmp_ln384_fu_128_p2;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_86;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_condition_86)) begin
        if (((icmp_ln373_fu_116_p2 == 1'd1) & (icmp_ln370_fu_104_p2 == 1'd0))) begin
            ap_phi_reg_pp0_iter1_p_Val2_s_reg_95 <= in_V_V_TDATA;
        end else if ((1'b1 == 1'b1)) begin
            ap_phi_reg_pp0_iter1_p_Val2_s_reg_95 <= ap_phi_reg_pp0_iter0_p_Val2_s_reg_95;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln370_fu_104_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        o_0_reg_73 <= select_ln384_fu_134_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        o_0_reg_73 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln370_reg_162 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        p_025_0_reg_61 <= {{ap_phi_mux_p_Val2_s_phi_fu_98_p4[15:8]}};
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        p_025_0_reg_61 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln370_fu_104_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        t_0_reg_84 <= t_fu_110_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        t_0_reg_84 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln370_reg_162 <= icmp_ln370_fu_104_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln370_fu_104_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln373_reg_171 <= icmp_ln373_fu_116_p2;
    end
end

always @ (*) begin
    if ((icmp_ln370_fu_104_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln373_reg_171 == 1'd0) & (icmp_ln370_reg_162 == 1'd0))) begin
        ap_phi_mux_p_Val2_s_phi_fu_98_p4 = zext_ln370_fu_142_p1;
    end else begin
        ap_phi_mux_p_Val2_s_phi_fu_98_p4 = ap_phi_reg_pp0_iter1_p_Val2_s_reg_95;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln373_fu_116_p2 == 1'd1) & (icmp_ln370_fu_104_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op16_read_state2 == 1'b1))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln370_reg_162 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln370_reg_162 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((icmp_ln370_fu_104_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((icmp_ln370_fu_104_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_op16_read_state2 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_op16_read_state2 == 1'b1)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_op16_read_state2 == 1'b1)));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = ((in_V_V_TVALID == 1'b0) & (ap_predicate_op16_read_state2 == 1'b1));
end

always @ (*) begin
    ap_block_state3_io = ((icmp_ln370_reg_162 == 1'd0) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_86 = ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_reg_pp0_iter0_p_Val2_s_reg_95 = 'bx;

always @ (*) begin
    ap_predicate_op16_read_state2 = ((icmp_ln373_fu_116_p2 == 1'd1) & (icmp_ln370_fu_104_p2 == 1'd0));
end

assign icmp_ln370_fu_104_p2 = ((t_0_reg_84 == 9'd256) ? 1'b1 : 1'b0);

assign icmp_ln373_fu_116_p2 = ((o_0_reg_73 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln384_fu_128_p2 = ((o_fu_122_p2 == 32'd2) ? 1'b1 : 1'b0);

assign o_fu_122_p2 = (32'd1 + o_0_reg_73);

assign out_V_V_TDATA = ap_phi_mux_p_Val2_s_phi_fu_98_p4[7:0];

assign select_ln384_fu_134_p3 = ((icmp_ln384_fu_128_p2[0:0] === 1'b1) ? 32'd0 : o_fu_122_p2);

assign t_fu_110_p2 = (t_0_reg_84 + 9'd1);

assign zext_ln370_fu_142_p1 = p_025_0_reg_61;

endmodule //StreamingDataWidthConverter_Batch_5_StreamingDataWidthCo_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcOgC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcOgC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcOgC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcOgC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcOgC_rom Thresholding_Batch_0_Thresholding_BatcOgC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActHfu.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActHfu_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActHfu_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActHfu(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActHfu_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActHfu_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActAem.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActAem_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActAem_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActAem(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActAem_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActAem_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_2_0/synth/finn_design_StreamingFCLayer_Batch_2_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFCLayer_Batch_3:1.0
// IP Revision: 2101301318

(* X_CORE_INFO = "StreamingFCLayer_Batch_3_StreamingFCLayer_Batch_3,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_2_0,StreamingFCLayer_Batch_3_StreamingFCLayer_Batch_3,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_2_0,StreamingFCLayer_Batch_3_StreamingFCLayer_Batch_3,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFCLayer_Batch_3,x_ipVersion=1.0,x_ipCoreRevision=2101301318,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_2_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  weights_V_V_TVALID,
  weights_V_V_TREADY,
  weights_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:weights_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 4, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [31 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TVALID" *)
input wire weights_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TREADY" *)
output wire weights_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME weights_V_V, TDATA_NUM_BYTES 16, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TDATA" *)
input wire [127 : 0] weights_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;

  StreamingFCLayer_Batch_3_StreamingFCLayer_Batch_3 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .weights_V_V_TVALID(weights_V_V_TVALID),
    .weights_V_V_TREADY(weights_V_V_TREADY),
    .weights_V_V_TDATA(weights_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActrcU.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActrcU_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActrcU_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActrcU(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActrcU_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActrcU_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbun.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbun_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbun_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbun(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbun_rom Thresholding_Batch_0_Thresholding_Batcbun_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Act0iy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Act0iy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Act0iy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Act0iy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Act0iy_rom StreamingFCLayer_Batch_4_Matrix_Vector_Act0iy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_BatcfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_BatcfYi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_BatcfYi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_BatcfYi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_BatcfYi_rom Thresholding_Batch_1_Thresholding_BatcfYi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActqcK.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActqcK_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActqcK_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActqcK(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActqcK_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActqcK_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_BatcjbC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_BatcjbC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_BatcjbC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_BatcjbC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_BatcjbC_rom Thresholding_Batch_2_Thresholding_BatcjbC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/e03c/hdl/verilog/ConvolutionInputGenerator_3_ConvolutionInputGenerator_3.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="ConvolutionInputGenerator_3_ConvolutionInputGenerator_3,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.054750,HLS_SYN_LAT=57173,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=606,HLS_SYN_LUT=1870,HLS_VERSION=2020_1_1}" *)

module ConvolutionInputGenerator_3_ConvolutionInputGenerator_3 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [31:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_ConvolutionInputGene_1_fu_26_ap_start;
wire    grp_ConvolutionInputGene_1_fu_26_ap_done;
wire    grp_ConvolutionInputGene_1_fu_26_ap_idle;
wire    grp_ConvolutionInputGene_1_fu_26_ap_ready;
wire    grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY;
wire   [31:0] grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA;
wire    grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID;
wire    grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY;
reg    grp_ConvolutionInputGene_1_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [31:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_ConvolutionInputGene_1_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

ConvolutionInputGenerator_3_ConvolutionInputGene_1 grp_ConvolutionInputGene_1_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_ConvolutionInputGene_1_fu_26_ap_start),
    .ap_done(grp_ConvolutionInputGene_1_fu_26_ap_done),
    .ap_idle(grp_ConvolutionInputGene_1_fu_26_ap_idle),
    .ap_ready(grp_ConvolutionInputGene_1_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 32 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 32 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA),
    .vld_in(grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_ConvolutionInputGene_1_fu_26_ap_ready == 1'b1)) begin
            grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_ConvolutionInputGene_1_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_ConvolutionInputGene_1_fu_26_ap_start = grp_ConvolutionInputGene_1_fu_26_ap_start_reg;

assign grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //ConvolutionInputGenerator_3_ConvolutionInputGenerator_3
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/5609/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccWB.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccWB_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccWB_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccWB(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccWB_rom Thresholding_Batch_0_Thresholding_BatccWB_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc7D.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcc7D_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc7D_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcc7D(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcc7D_rom Thresholding_Batch_0_Thresholding_Batcc7D_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actibs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actibs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actibs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actibs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actibs_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actibs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_6_wstrm_0/synth/finn_design_StreamingFCLayer_Batch_6_wstrm_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:user:memstream:1.0
// IP Revision: 5

(* X_CORE_INFO = "memstream,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_6_wstrm_0,memstream,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_6_wstrm_0,memstream,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=user,x_ipName=memstream,x_ipVersion=1.0,x_ipCoreRevision=5,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED,CONFIG_EN=true,NSTREAMS=1,MEM_DEPTH=1792,MEM_WIDTH=8,MEM_INIT=/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_6_e2ail04f/,RAM_STYLE=distributed,STRM0_WIDTH=8,STRM1_WIDTH=32,STRM2_WIDTH=32,STRM3_WIDTH=32,STRM4_WIDTH=32,STRM5_WIDTH=32\
,STRM0_DEPTH=1792,STRM1_DEPTH=2304,STRM2_DEPTH=2304,STRM3_DEPTH=2304,STRM4_DEPTH=2304,STRM5_DEPTH=2304,STRM0_OFFSET=0,STRM1_OFFSET=2304,STRM2_OFFSET=4608,STRM3_OFFSET=6912,STRM4_OFFSET=9216,STRM5_OFFSET=11520,AXILITE_ADDR_WIDTH=13}" *)
(* IP_DEFINITION_SOURCE = "package_project" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_6_wstrm_0 (
  aclk,
  aresetn,
  awready,
  awvalid,
  awaddr,
  awprot,
  wready,
  wvalid,
  wdata,
  wstrb,
  bready,
  bvalid,
  bresp,
  arready,
  arvalid,
  araddr,
  arprot,
  rready,
  rvalid,
  rresp,
  rdata,
  m_axis_0_tready,
  m_axis_0_tvalid,
  m_axis_0_tdata
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aclk, ASSOCIATED_BUSIF m_axis_0:m_axis_1:m_axis_2:m_axis_3:m_axis_4:m_axis_5:s_axilite, ASSOCIATED_RESET aresetn, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 aclk CLK" *)
input wire aclk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aresetn, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 aresetn RST" *)
input wire aresetn;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWREADY" *)
output wire awready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWVALID" *)
input wire awvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWADDR" *)
input wire [12 : 0] awaddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWPROT" *)
input wire [2 : 0] awprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WREADY" *)
output wire wready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WVALID" *)
input wire wvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WDATA" *)
input wire [31 : 0] wdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WSTRB" *)
input wire [3 : 0] wstrb;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BREADY" *)
input wire bready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BVALID" *)
output wire bvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BRESP" *)
output wire [1 : 0] bresp;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARREADY" *)
output wire arready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARVALID" *)
input wire arvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARADDR" *)
input wire [12 : 0] araddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARPROT" *)
input wire [2 : 0] arprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RREADY" *)
input wire rready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RVALID" *)
output wire rvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RRESP" *)
output wire [1 : 0] rresp;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axilite, DATA_WIDTH 32, PROTOCOL AXI4LITE, FREQ_HZ 100000000.000000, ID_WIDTH 0, ADDR_WIDTH 13, AWUSER_WIDTH 0, ARUSER_WIDTH 0, WUSER_WIDTH 0, RUSER_WIDTH 0, BUSER_WIDTH 0, READ_WRITE_MODE READ_WRITE, HAS_BURST 0, HAS_LOCK 0, HAS_PROT 1, HAS_CACHE 0, HAS_QOS 0, HAS_REGION 0, HAS_WSTRB 1, HAS_BRESP 1, HAS_RRESP 1, SUPPORTS_NARROW_BURST 0, NUM_READ_OUTSTANDING 1, NUM_WRITE_OUTSTANDING 1, MAX_BURST_LENGTH 1, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, NUM_READ_THREADS 1, NUM_W\
RITE_THREADS 1, RUSER_BITS_PER_BYTE 0, WUSER_BITS_PER_BYTE 0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RDATA" *)
output wire [31 : 0] rdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TREADY" *)
input wire m_axis_0_tready;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TVALID" *)
output wire m_axis_0_tvalid;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME m_axis_0, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TDATA" *)
output wire [7 : 0] m_axis_0_tdata;

  memstream #(
    .CONFIG_EN(1'B1),
    .NSTREAMS(1),
    .MEM_DEPTH(1792),
    .MEM_WIDTH(8),
    .MEM_INIT("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_6_e2ail04f/"),
    .RAM_STYLE("distributed"),
    .STRM0_WIDTH(8),
    .STRM1_WIDTH(32),
    .STRM2_WIDTH(32),
    .STRM3_WIDTH(32),
    .STRM4_WIDTH(32),
    .STRM5_WIDTH(32),
    .STRM0_DEPTH(1792),
    .STRM1_DEPTH(2304),
    .STRM2_DEPTH(2304),
    .STRM3_DEPTH(2304),
    .STRM4_DEPTH(2304),
    .STRM5_DEPTH(2304),
    .STRM0_OFFSET(0),
    .STRM1_OFFSET(2304),
    .STRM2_OFFSET(4608),
    .STRM3_OFFSET(6912),
    .STRM4_OFFSET(9216),
    .STRM5_OFFSET(11520),
    .AXILITE_ADDR_WIDTH(13)
  ) inst (
    .aclk(aclk),
    .aresetn(aresetn),
    .awready(awready),
    .awvalid(awvalid),
    .awaddr(awaddr),
    .awprot(awprot),
    .wready(wready),
    .wvalid(wvalid),
    .wdata(wdata),
    .wstrb(wstrb),
    .bready(bready),
    .bvalid(bvalid),
    .bresp(bresp),
    .arready(arready),
    .arvalid(arvalid),
    .araddr(araddr),
    .arprot(arprot),
    .rready(rready),
    .rvalid(rvalid),
    .rresp(rresp),
    .rdata(rdata),
    .m_axis_0_afull(1'B0),
    .m_axis_0_tready(m_axis_0_tready),
    .m_axis_0_tvalid(m_axis_0_tvalid),
    .m_axis_0_tdata(m_axis_0_tdata),
    .m_axis_1_afull(1'B0),
    .m_axis_1_tready(1'B1),
    .m_axis_1_tvalid(),
    .m_axis_1_tdata(),
    .m_axis_2_afull(1'B0),
    .m_axis_2_tready(1'B1),
    .m_axis_2_tvalid(),
    .m_axis_2_tdata(),
    .m_axis_3_afull(1'B0),
    .m_axis_3_tready(1'B1),
    .m_axis_3_tvalid(),
    .m_axis_3_tdata(),
    .m_axis_4_afull(1'B0),
    .m_axis_4_tready(1'B1),
    .m_axis_4_tvalid(),
    .m_axis_4_tdata(),
    .m_axis_5_afull(1'B0),
    .m_axis_5_tready(1'B1),
    .m_axis_5_tvalid(),
    .m_axis_5_tdata()
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actmb6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actmb6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actmb6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actmb6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actmb6_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actmb6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_19_0/synth/finn_design_StreamingFIFO_19_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_19:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_19,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_19_0,StreamingFIFO_19,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_19_0,StreamingFIFO_19,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_19,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_19_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [7 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_19 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccMA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccMA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccMA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccMA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccMA_rom Thresholding_Batch_0_Thresholding_BatccMA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActHfu.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActHfu_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActHfu_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActHfu(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActHfu_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActHfu_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_11_0/synth/finn_design_StreamingFIFO_11_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_11:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_11,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_11_0,StreamingFIFO_11,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_11_0,StreamingFIFO_11,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_11,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_11_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_11 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/eb12/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actg8j.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actg8j_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actg8j_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actg8j(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actg8j_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actg8j_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActRg6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActRg6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActRg6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActRg6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActRg6_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActRg6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/e03c/hdl/verilog/ConvolutionInputGenerator_3_ConvolutionInputGfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module ConvolutionInputGenerator_3_ConvolutionInputGfYi #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [31 : 0]     din0,
    input  [31 : 0]     din1,
    input  [31 : 0]     din2,
    input  [31 : 0]     din3,
    input  [1 : 0]    din4,
    output [31 : 0]   dout);

// puts internal signals
wire [1 : 0]     sel;
// level 1 signals
wire [31 : 0]         mux_1_0;
wire [31 : 0]         mux_1_1;
// level 2 signals
wire [31 : 0]         mux_2_0;

assign sel = din4;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;

// output logic
assign dout = mux_2_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/6405/hdl/verilog/StreamingFCLayer_Batch_5_StreamingFCLayer_Batch_5.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingFCLayer_Batch_5_StreamingFCLayer_Batch_5,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.042250,HLS_SYN_LAT=3612678,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=2520,HLS_SYN_LUT=1083,HLS_VERSION=2020_1_1}" *)

module StreamingFCLayer_Batch_5_StreamingFCLayer_Batch_5 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        weights_V_V_TDATA,
        weights_V_V_TVALID,
        weights_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [31:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
input  [31:0] weights_V_V_TDATA;
input   weights_V_V_TVALID;
output   weights_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;
reg weights_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_Matrix_Vector_Activa_fu_28_ap_start;
wire    grp_Matrix_Vector_Activa_fu_28_ap_done;
wire    grp_Matrix_Vector_Activa_fu_28_ap_idle;
wire    grp_Matrix_Vector_Activa_fu_28_ap_ready;
wire    grp_Matrix_Vector_Activa_fu_28_in_V_V_TREADY;
wire   [15:0] grp_Matrix_Vector_Activa_fu_28_out_V_V_TDATA;
wire    grp_Matrix_Vector_Activa_fu_28_out_V_V_TVALID;
wire    grp_Matrix_Vector_Activa_fu_28_out_V_V_TREADY;
wire    grp_Matrix_Vector_Activa_fu_28_weight_V_V_TREADY;
reg    grp_Matrix_Vector_Activa_fu_28_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [31:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    regslice_both_weights_V_V_U_apdone_blk;
wire   [31:0] weights_V_V_TDATA_int;
wire    weights_V_V_TVALID_int;
reg    weights_V_V_TREADY_int;
wire    regslice_both_weights_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_Matrix_Vector_Activa_fu_28_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingFCLayer_Batch_5_Matrix_Vector_Activa grp_Matrix_Vector_Activa_fu_28(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_Matrix_Vector_Activa_fu_28_ap_start),
    .ap_done(grp_Matrix_Vector_Activa_fu_28_ap_done),
    .ap_idle(grp_Matrix_Vector_Activa_fu_28_ap_idle),
    .ap_ready(grp_Matrix_Vector_Activa_fu_28_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_Matrix_Vector_Activa_fu_28_in_V_V_TREADY),
    .out_V_V_TDATA(grp_Matrix_Vector_Activa_fu_28_out_V_V_TDATA),
    .out_V_V_TVALID(grp_Matrix_Vector_Activa_fu_28_out_V_V_TVALID),
    .out_V_V_TREADY(grp_Matrix_Vector_Activa_fu_28_out_V_V_TREADY),
    .weight_V_V_TDATA(weights_V_V_TDATA_int),
    .weight_V_V_TVALID(weights_V_V_TVALID_int),
    .weight_V_V_TREADY(grp_Matrix_Vector_Activa_fu_28_weight_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 32 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 32 ))
regslice_both_weights_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(weights_V_V_TDATA),
    .vld_in(weights_V_V_TVALID),
    .ack_in(regslice_both_weights_V_V_U_ack_in),
    .data_out(weights_V_V_TDATA_int),
    .vld_out(weights_V_V_TVALID_int),
    .ack_out(weights_V_V_TREADY_int),
    .apdone_blk(regslice_both_weights_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_Matrix_Vector_Activa_fu_28_out_V_V_TDATA),
    .vld_in(grp_Matrix_Vector_Activa_fu_28_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_Matrix_Vector_Activa_fu_28_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_Matrix_Vector_Activa_fu_28_ap_start_reg <= 1'b1;
        end else if ((grp_Matrix_Vector_Activa_fu_28_ap_ready == 1'b1)) begin
            grp_Matrix_Vector_Activa_fu_28_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_28_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    if (((regslice_both_weights_V_V_U_ack_in == 1'b1) & (weights_V_V_TVALID == 1'b1))) begin
        weights_V_V_TREADY = 1'b1;
    end else begin
        weights_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        weights_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_28_weight_V_V_TREADY;
    end else begin
        weights_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_Matrix_Vector_Activa_fu_28_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_Matrix_Vector_Activa_fu_28_ap_start = grp_Matrix_Vector_Activa_fu_28_ap_start_reg;

assign grp_Matrix_Vector_Activa_fu_28_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingFCLayer_Batch_5_StreamingFCLayer_Batch_5
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActdEe.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActdEe_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActdEe_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActdEe(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActdEe_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActdEe_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcIfE.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcIfE_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcIfE_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcIfE(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcIfE_rom Thresholding_Batch_0_Thresholding_BatcIfE_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Acttde.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Acttde_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Acttde_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Acttde(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Acttde_rom StreamingFCLayer_Batch_3_Matrix_Vector_Acttde_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Act1iI.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Act1iI_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Act1iI_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Act1iI(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Act1iI_rom StreamingFCLayer_Batch_2_Matrix_Vector_Act1iI_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/841a/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActUhA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActUhA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActUhA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActUhA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActUhA_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActUhA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcMgi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcMgi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcMgi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcMgi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcMgi_rom Thresholding_Batch_0_Thresholding_BatcMgi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_BatcdEe.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_BatcdEe_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_BatcdEe_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_BatcdEe(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_BatcdEe_rom Thresholding_Batch_1_Thresholding_BatcdEe_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccyx.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccyx_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccyx_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccyx(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccyx_rom Thresholding_Batch_0_Thresholding_Batccyx_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActeOg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActeOg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActeOg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActeOg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActeOg_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActeOg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActAem.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActAem_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActAem_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActAem(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActAem_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActAem_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActYie.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActYie_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActYie_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActYie(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActYie_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActYie_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actmb6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actmb6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actmb6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actmb6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actmb6_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actmb6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcmb6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_Batcmb6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcmb6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_Batcmb6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_Batcmb6_rom Thresholding_Batch_2_Thresholding_Batcmb6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccFz.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccFz_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccFz_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccFz(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccFz_rom Thresholding_Batch_0_Thresholding_BatccFz_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/f5c4/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_BatcjbC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_BatcjbC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_BatcjbC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_BatcjbC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_BatcjbC_rom Thresholding_Batch_1_Thresholding_BatcjbC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/c3f7/hdl/verilog/LabelSelect_Batch_0_LabelSelect_Batch_0.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="LabelSelect_Batch_0_LabelSelect_Batch_0,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=3.677000,HLS_SYN_LAT=12,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=35,HLS_SYN_LUT=155,HLS_VERSION=2020_1_1}" *)

module LabelSelect_Batch_0_LabelSelect_Batch_0 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_LabelSelect_Batch_fu_26_ap_start;
wire    grp_LabelSelect_Batch_fu_26_ap_done;
wire    grp_LabelSelect_Batch_fu_26_ap_idle;
wire    grp_LabelSelect_Batch_fu_26_ap_ready;
wire    grp_LabelSelect_Batch_fu_26_in_V_V_TREADY;
wire   [7:0] grp_LabelSelect_Batch_fu_26_out_V_V_TDATA;
wire    grp_LabelSelect_Batch_fu_26_out_V_V_TVALID;
wire    grp_LabelSelect_Batch_fu_26_out_V_V_TREADY;
reg    grp_LabelSelect_Batch_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [15:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_LabelSelect_Batch_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

LabelSelect_Batch_0_LabelSelect_Batch grp_LabelSelect_Batch_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_LabelSelect_Batch_fu_26_ap_start),
    .ap_done(grp_LabelSelect_Batch_fu_26_ap_done),
    .ap_idle(grp_LabelSelect_Batch_fu_26_ap_idle),
    .ap_ready(grp_LabelSelect_Batch_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_LabelSelect_Batch_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_LabelSelect_Batch_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_LabelSelect_Batch_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_LabelSelect_Batch_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_LabelSelect_Batch_fu_26_out_V_V_TDATA),
    .vld_in(grp_LabelSelect_Batch_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_LabelSelect_Batch_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_LabelSelect_Batch_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_LabelSelect_Batch_fu_26_ap_ready == 1'b1)) begin
            grp_LabelSelect_Batch_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_LabelSelect_Batch_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_LabelSelect_Batch_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_LabelSelect_Batch_fu_26_ap_start = grp_LabelSelect_Batch_fu_26_ap_start_reg;

assign grp_LabelSelect_Batch_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //LabelSelect_Batch_0_LabelSelect_Batch_0
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccOA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccOA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccOA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccOA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccOA_rom Thresholding_Batch_0_Thresholding_BatccOA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActkbM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActkbM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActkbM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActkbM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActkbM_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActkbM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActKfY.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActKfY_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActKfY_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActKfY(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActKfY_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActKfY_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_6_0/synth/finn_design_StreamingFIFO_6_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_6:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_6,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_6_0,StreamingFIFO_6,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_6_0,StreamingFIFO_6,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_6,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_6_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [23 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 3, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [23 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 3, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_6 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActVhK.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActVhK_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActVhK_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActVhK(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActVhK_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActVhK_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActrcU.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActrcU_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActrcU_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActrcU(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActrcU_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActrcU_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdfE.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcdfE_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcdfE_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcdfE(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcdfE_rom Thresholding_Batch_0_Thresholding_BatcdfE_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcPgM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcPgM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcPgM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcPgM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcPgM_rom Thresholding_Batch_0_Thresholding_BatcPgM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Act3i2.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Act3i2_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Act3i2_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Act3i2(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Act3i2_rom StreamingFCLayer_Batch_1_Matrix_Vector_Act3i2_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingDataWidthConverter_Batch_3_0/synth/finn_design_StreamingDataWidthConverter_Batch_3_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingDataWidthConverter_Batch_3:1.0
// IP Revision: 2101301321

(* X_CORE_INFO = "StreamingDataWidthConverter_Batch_3_StreamingDataWidthConverter_Batch_3,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingDataWidthConverter_Batch_3_0,StreamingDataWidthConverter_Batch_3_StreamingDataWidthConverter_Batch_3,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingDataWidthConverter_Batch_3_0,StreamingDataWidthConverter_Batch_3_StreamingDataWidthConverter_Batch_3,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingDataWidthConverter_Batch_3,x_ipVersion=1.0,x_ipCoreRevision=2101301321,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingDataWidthConverter_Batch_3_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 4, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [31 : 0] out_V_V_TDATA;

  StreamingDataWidthConverter_Batch_3_StreamingDataWidthConverter_Batch_3 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActYie.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActYie_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActYie_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActYie(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActYie_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActYie_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccAy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccAy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccAy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccAy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccAy_rom Thresholding_Batch_0_Thresholding_BatccAy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingDataWidthConverter_Batch_1_0/synth/finn_design_StreamingDataWidthConverter_Batch_1_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingDataWidthConverter_Batch_1:1.0
// IP Revision: 2101301322

(* X_CORE_INFO = "StreamingDataWidthConverter_Batch_1_StreamingDataWidthConverter_Batch_1,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingDataWidthConverter_Batch_1_0,StreamingDataWidthConverter_Batch_1_StreamingDataWidthConverter_Batch_1,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingDataWidthConverter_Batch_1_0,StreamingDataWidthConverter_Batch_1_StreamingDataWidthConverter_Batch_1,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingDataWidthConverter_Batch_1,x_ipVersion=1.0,x_ipCoreRevision=2101301322,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingDataWidthConverter_Batch_1_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 12, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [95 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 3, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [23 : 0] out_V_V_TDATA;

  StreamingDataWidthConverter_Batch_1_StreamingDataWidthConverter_Batch_1 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActVhK.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActVhK_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActVhK_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActVhK(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActVhK_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActVhK_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActfYi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActfYi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActfYi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActfYi_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActfYi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActDeQ.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActDeQ_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActDeQ_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActDeQ(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActDeQ_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActDeQ_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActPgM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActPgM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActPgM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActPgM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActPgM_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActPgM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccSB.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccSB_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccSB_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccSB(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccSB_rom Thresholding_Batch_0_Thresholding_BatccSB_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccow.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccow_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccow_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccow(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccow_rom Thresholding_Batch_0_Thresholding_Batccow_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_4_0/synth/finn_design_StreamingFIFO_4_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_4:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_4,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_4_0,StreamingFIFO_4,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_4_0,StreamingFIFO_4,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_4,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_4_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [95 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 12, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [95 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 12, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_4 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_BatceOg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_BatceOg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_BatceOg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_BatceOg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_BatceOg_rom Thresholding_Batch_1_Thresholding_BatceOg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_5_0/synth/finn_design_StreamingFIFO_5_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_5:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_5,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_5_0,StreamingFIFO_5,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_5_0,StreamingFIFO_5,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_5,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_5_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_5 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actmb6.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actmb6_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actmb6_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actmb6(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actmb6_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actmb6_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/abe7/hdl/verilog/ConvolutionInputGenerator_0_ConvolutionInputGfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module ConvolutionInputGenerator_0_ConvolutionInputGfYi #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [7 : 0]     din0,
    input  [7 : 0]     din1,
    input  [7 : 0]     din2,
    input  [7 : 0]     din3,
    input  [1 : 0]    din4,
    output [7 : 0]   dout);

// puts internal signals
wire [1 : 0]     sel;
// level 1 signals
wire [7 : 0]         mux_1_0;
wire [7 : 0]         mux_1_1;
// level 2 signals
wire [7 : 0]         mux_2_0;

assign sel = din4;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;

// output logic
assign dout = mux_2_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcKfY.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcKfY_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcKfY_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcKfY(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcKfY_rom Thresholding_Batch_0_Thresholding_BatcKfY_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actcud.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actcud_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actcud_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actcud(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actcud_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actcud_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbom.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbom_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbom_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbom(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbom_rom Thresholding_Batch_0_Thresholding_Batcbom_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/2539/hdl/verilog/StreamingDataWidthConverter_Batch_4_StreamingDataWidthCo_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingDataWidthConverter_Batch_4_StreamingDataWidthCo_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [15:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln402_fu_88_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln411_reg_154;
reg   [15:0] r_V_reg_61;
reg   [13:0] t_0_reg_72;
reg   [0:0] icmp_ln402_reg_135;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [13:0] t_fu_94_p2;
reg   [15:0] tmp_V_reg_144;
wire   [31:0] p_Result_s_fu_103_p3;
reg   [31:0] p_Result_s_reg_149;
wire   [0:0] icmp_ln411_fu_117_p2;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg   [15:0] ap_phi_mux_r_V_phi_fu_65_p4;
reg   [31:0] i_1_fu_44;
wire   [31:0] i_fu_111_p2;
reg    ap_block_pp0_stage0_01001;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_fu_117_p2 == 1'd0) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_1_fu_44 <= i_fu_111_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_fu_117_p2 == 1'd1) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        i_1_fu_44 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_reg_135 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        r_V_reg_61 <= tmp_V_reg_144;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        r_V_reg_61 <= 16'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        t_0_reg_72 <= t_fu_94_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        t_0_reg_72 <= 14'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln402_reg_135 <= icmp_ln402_fu_88_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln411_reg_154 <= icmp_ln411_fu_117_p2;
        p_Result_s_reg_149 <= p_Result_s_fu_103_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_reg_144 <= in_V_V_TDATA;
    end
end

always @ (*) begin
    if ((icmp_ln402_fu_88_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln402_reg_135 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_r_V_phi_fu_65_p4 = tmp_V_reg_144;
    end else begin
        ap_phi_mux_r_V_phi_fu_65_p4 = r_V_reg_61;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln402_fu_88_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln402_fu_88_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln411_reg_154 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln411_reg_154 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln402_fu_88_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln402_fu_88_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = ((icmp_ln402_fu_88_p2 == 1'd0) & (in_V_V_TVALID == 1'b0));
end

always @ (*) begin
    ap_block_state3_io = ((icmp_ln411_reg_154 == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign i_fu_111_p2 = (i_1_fu_44 + 32'd1);

assign icmp_ln402_fu_88_p2 = ((t_0_reg_72 == 14'd14400) ? 1'b1 : 1'b0);

assign icmp_ln411_fu_117_p2 = ((i_fu_111_p2 == 32'd2) ? 1'b1 : 1'b0);

assign out_V_V_TDATA = p_Result_s_reg_149;

assign p_Result_s_fu_103_p3 = {{in_V_V_TDATA}, {ap_phi_mux_r_V_phi_fu_65_p4}};

assign t_fu_94_p2 = (t_0_reg_72 + 14'd1);

endmodule //StreamingDataWidthConverter_Batch_4_StreamingDataWidthCo_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_5_0/synth/finn_design_StreamingFCLayer_Batch_5_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFCLayer_Batch_5:1.0
// IP Revision: 2101301315

(* X_CORE_INFO = "StreamingFCLayer_Batch_5_StreamingFCLayer_Batch_5,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_5_0,StreamingFCLayer_Batch_5_StreamingFCLayer_Batch_5,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_5_0,StreamingFCLayer_Batch_5_StreamingFCLayer_Batch_5,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFCLayer_Batch_5,x_ipVersion=1.0,x_ipCoreRevision=2101301315,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_5_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  weights_V_V_TVALID,
  weights_V_V_TREADY,
  weights_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:weights_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 4, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [31 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TVALID" *)
input wire weights_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TREADY" *)
output wire weights_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME weights_V_V, TDATA_NUM_BYTES 4, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 weights_V_V TDATA" *)
input wire [31 : 0] weights_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;

  StreamingFCLayer_Batch_5_StreamingFCLayer_Batch_5 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .weights_V_V_TVALID(weights_V_V_TVALID),
    .weights_V_V_TREADY(weights_V_V_TREADY),
    .weights_V_V_TDATA(weights_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_Batccud.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_Batccud_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_Batccud_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_Batccud(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_Batccud_rom Thresholding_Batch_2_Thresholding_Batccud_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/2539/hdl/verilog/StreamingDataWidthConverter_Batch_4_StreamingDataWidthConverter_Batch_4.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingDataWidthConverter_Batch_4_StreamingDataWidthConverter_Batch_4,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=5.025000,HLS_SYN_LAT=14405,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=122,HLS_SYN_LUT=229,HLS_VERSION=2020_1_1}" *)

module StreamingDataWidthConverter_Batch_4_StreamingDataWidthConverter_Batch_4 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_start;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_done;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_idle;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_ready;
wire    grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
wire   [31:0] grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY;
reg    grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [15:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_StreamingDataWidthCo_1_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingDataWidthConverter_Batch_4_StreamingDataWidthCo_1 grp_StreamingDataWidthCo_1_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_StreamingDataWidthCo_1_fu_26_ap_start),
    .ap_done(grp_StreamingDataWidthCo_1_fu_26_ap_done),
    .ap_idle(grp_StreamingDataWidthCo_1_fu_26_ap_idle),
    .ap_ready(grp_StreamingDataWidthCo_1_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 32 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .vld_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_StreamingDataWidthCo_1_fu_26_ap_ready == 1'b1)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_StreamingDataWidthCo_1_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_StreamingDataWidthCo_1_fu_26_ap_start = grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;

assign grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingDataWidthConverter_Batch_4_StreamingDataWidthConverter_Batch_4
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/466a/hdl/verilog/StreamingDataWidthConverter_Batch_1_StreamingDataWidthConverter_Batch_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingDataWidthConverter_Batch_1_StreamingDataWidthConverter_Batch_1,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=5.723000,HLS_SYN_LAT=12805,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=226,HLS_SYN_LUT=292,HLS_VERSION=2020_1_1}" *)

module StreamingDataWidthConverter_Batch_1_StreamingDataWidthConverter_Batch_1 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [95:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [23:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_start;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_done;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_idle;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_ready;
wire    grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
wire   [23:0] grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY;
reg    grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [95:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_StreamingDataWidthCo_1_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingDataWidthConverter_Batch_1_StreamingDataWidthCo_1 grp_StreamingDataWidthCo_1_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_StreamingDataWidthCo_1_fu_26_ap_start),
    .ap_done(grp_StreamingDataWidthCo_1_fu_26_ap_done),
    .ap_idle(grp_StreamingDataWidthCo_1_fu_26_ap_idle),
    .ap_ready(grp_StreamingDataWidthCo_1_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 96 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 24 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .vld_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_StreamingDataWidthCo_1_fu_26_ap_ready == 1'b1)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_StreamingDataWidthCo_1_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_StreamingDataWidthCo_1_fu_26_ap_start = grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;

assign grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingDataWidthConverter_Batch_1_StreamingDataWidthConverter_Batch_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActGfk.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActGfk_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActGfk_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActGfk(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActGfk_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActGfk_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcQgW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcQgW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcQgW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcQgW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcQgW_rom Thresholding_Batch_0_Thresholding_BatcQgW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActGfk.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActGfk_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActGfk_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActGfk(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActGfk_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActGfk_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8ee6/StreamingFIFO_10.v


module StreamingFIFO_10(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(16)
)
StreamingFIFO_10_StreamingFIFO_10
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActNgs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActNgs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActNgs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActNgs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActNgs_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActNgs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcGfk.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcGfk_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcGfk_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcGfk(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcGfk_rom Thresholding_Batch_0_Thresholding_BatcGfk_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/2c22/hdl/verilog/ConvolutionInputGenerator_2_ConvolutionInputGbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module ConvolutionInputGenerator_2_ConvolutionInputGbkb_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 24;
parameter AWIDTH = 5;
parameter MEM_SIZE = 32;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];




always @(posedge clk)  
begin 
    if (ce0) begin
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module ConvolutionInputGenerator_2_ConvolutionInputGbkb(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd24;
parameter AddressRange = 32'd32;
parameter AddressWidth = 32'd5;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



ConvolutionInputGenerator_2_ConvolutionInputGbkb_ram ConvolutionInputGenerator_2_ConvolutionInputGbkb_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActrcU.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActrcU_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActrcU_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActrcU(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActrcU_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActrcU_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_BatcdEe.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_BatcdEe_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_BatcdEe_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_BatcdEe(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_BatcdEe_rom Thresholding_Batch_2_Thresholding_BatcdEe_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Act1iI.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Act1iI_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Act1iI_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Act1iI(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Act1iI_rom StreamingFCLayer_Batch_3_Matrix_Vector_Act1iI_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_2_0/synth/finn_design_StreamingFIFO_2_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_2:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_2,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_2_0,StreamingFIFO_2,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_2_0,StreamingFIFO_2,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_2,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_2_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [15 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [15 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_2 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/46bc/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcctx.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcctx_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcctx_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcctx(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcctx_rom Thresholding_Batch_0_Thresholding_Batcctx_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/1ba7/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccHz.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccHz_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccHz_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccHz(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccHz_rom Thresholding_Batch_0_Thresholding_BatccHz_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActYie.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActYie_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActYie_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActYie(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActYie_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActYie_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/abe7/hdl/verilog/ConvolutionInputGenerator_0_ConvolutionInputGbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module ConvolutionInputGenerator_0_ConvolutionInputGbkb_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 8;
parameter AWIDTH = 10;
parameter MEM_SIZE = 768;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];




always @(posedge clk)  
begin 
    if (ce0) begin
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module ConvolutionInputGenerator_0_ConvolutionInputGbkb(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd768;
parameter AddressWidth = 32'd10;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



ConvolutionInputGenerator_0_ConvolutionInputGbkb_ram ConvolutionInputGenerator_0_ConvolutionInputGbkb_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/cd9c/hdl/verilog/StreamingFCLayer_Batch_0_StreamingFCLayer_Batch_0.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingFCLayer_Batch_0_StreamingFCLayer_Batch_0,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.573500,HLS_SYN_LAT=1843205,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=4841,HLS_SYN_LUT=3568,HLS_VERSION=2020_1_1}" *)

module StreamingFCLayer_Batch_0_StreamingFCLayer_Batch_0 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        weights_V_V_TDATA,
        weights_V_V_TVALID,
        weights_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [7:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
input  [31:0] weights_V_V_TDATA;
input   weights_V_V_TVALID;
output   weights_V_V_TREADY;
output  [95:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;
reg weights_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_Matrix_Vector_Activa_fu_28_ap_start;
wire    grp_Matrix_Vector_Activa_fu_28_ap_done;
wire    grp_Matrix_Vector_Activa_fu_28_ap_idle;
wire    grp_Matrix_Vector_Activa_fu_28_ap_ready;
wire    grp_Matrix_Vector_Activa_fu_28_in_V_V_TREADY;
wire   [95:0] grp_Matrix_Vector_Activa_fu_28_out_V_V_TDATA;
wire    grp_Matrix_Vector_Activa_fu_28_out_V_V_TVALID;
wire    grp_Matrix_Vector_Activa_fu_28_out_V_V_TREADY;
wire    grp_Matrix_Vector_Activa_fu_28_weight_V_V_TREADY;
reg    grp_Matrix_Vector_Activa_fu_28_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [7:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    regslice_both_weights_V_V_U_apdone_blk;
wire   [31:0] weights_V_V_TDATA_int;
wire    weights_V_V_TVALID_int;
reg    weights_V_V_TREADY_int;
wire    regslice_both_weights_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_Matrix_Vector_Activa_fu_28_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingFCLayer_Batch_0_Matrix_Vector_Activa grp_Matrix_Vector_Activa_fu_28(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_Matrix_Vector_Activa_fu_28_ap_start),
    .ap_done(grp_Matrix_Vector_Activa_fu_28_ap_done),
    .ap_idle(grp_Matrix_Vector_Activa_fu_28_ap_idle),
    .ap_ready(grp_Matrix_Vector_Activa_fu_28_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_Matrix_Vector_Activa_fu_28_in_V_V_TREADY),
    .out_V_V_TDATA(grp_Matrix_Vector_Activa_fu_28_out_V_V_TDATA),
    .out_V_V_TVALID(grp_Matrix_Vector_Activa_fu_28_out_V_V_TVALID),
    .out_V_V_TREADY(grp_Matrix_Vector_Activa_fu_28_out_V_V_TREADY),
    .weight_V_V_TDATA(weights_V_V_TDATA_int),
    .weight_V_V_TVALID(weights_V_V_TVALID_int),
    .weight_V_V_TREADY(grp_Matrix_Vector_Activa_fu_28_weight_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 8 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 32 ))
regslice_both_weights_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(weights_V_V_TDATA),
    .vld_in(weights_V_V_TVALID),
    .ack_in(regslice_both_weights_V_V_U_ack_in),
    .data_out(weights_V_V_TDATA_int),
    .vld_out(weights_V_V_TVALID_int),
    .ack_out(weights_V_V_TREADY_int),
    .apdone_blk(regslice_both_weights_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 96 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_Matrix_Vector_Activa_fu_28_out_V_V_TDATA),
    .vld_in(grp_Matrix_Vector_Activa_fu_28_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_Matrix_Vector_Activa_fu_28_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_Matrix_Vector_Activa_fu_28_ap_start_reg <= 1'b1;
        end else if ((grp_Matrix_Vector_Activa_fu_28_ap_ready == 1'b1)) begin
            grp_Matrix_Vector_Activa_fu_28_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_28_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    if (((regslice_both_weights_V_V_U_ack_in == 1'b1) & (weights_V_V_TVALID == 1'b1))) begin
        weights_V_V_TREADY = 1'b1;
    end else begin
        weights_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        weights_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_28_weight_V_V_TREADY;
    end else begin
        weights_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_Matrix_Vector_Activa_fu_28_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_Matrix_Vector_Activa_fu_28_ap_start = grp_Matrix_Vector_Activa_fu_28_ap_start_reg;

assign grp_Matrix_Vector_Activa_fu_28_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingFCLayer_Batch_0_StreamingFCLayer_Batch_0
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_StreamingFCLayer_6jw.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

(* use_dsp = "no" *) module StreamingFCLayer_Batch_3_StreamingFCLayer_6jw_Mul_LUT_0(a, b, p);
input[4 - 1 : 0] a; 
input[4 - 1 : 0] b; 
output[8 - 1 : 0] p;

assign p = $signed({1'b0, a}) * $signed(b);
endmodule
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_StreamingFCLayer_6jw(
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



StreamingFCLayer_Batch_3_StreamingFCLayer_6jw_Mul_LUT_0 StreamingFCLayer_Batch_3_StreamingFCLayer_6jw_Mul_LUT_0_U(
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFCLayer_Batch_2_wstrm_0/synth/finn_design_StreamingFCLayer_Batch_2_wstrm_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:user:memstream:1.0
// IP Revision: 5

(* X_CORE_INFO = "memstream,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFCLayer_Batch_2_wstrm_0,memstream,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFCLayer_Batch_2_wstrm_0,memstream,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=user,x_ipName=memstream,x_ipVersion=1.0,x_ipCoreRevision=5,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED,CONFIG_EN=true,NSTREAMS=1,MEM_DEPTH=4096,MEM_WIDTH=128,MEM_INIT=/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/,RAM_STYLE=block,STRM0_WIDTH=128,STRM1_WIDTH=32,STRM2_WIDTH=32,STRM3_WIDTH=32,STRM4_WIDTH=32,STRM5_WIDTH=32,S\
TRM0_DEPTH=4096,STRM1_DEPTH=2304,STRM2_DEPTH=2304,STRM3_DEPTH=2304,STRM4_DEPTH=2304,STRM5_DEPTH=2304,STRM0_OFFSET=0,STRM1_OFFSET=2304,STRM2_OFFSET=4608,STRM3_OFFSET=6912,STRM4_OFFSET=9216,STRM5_OFFSET=11520,AXILITE_ADDR_WIDTH=16}" *)
(* IP_DEFINITION_SOURCE = "package_project" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFCLayer_Batch_2_wstrm_0 (
  aclk,
  aresetn,
  awready,
  awvalid,
  awaddr,
  awprot,
  wready,
  wvalid,
  wdata,
  wstrb,
  bready,
  bvalid,
  bresp,
  arready,
  arvalid,
  araddr,
  arprot,
  rready,
  rvalid,
  rresp,
  rdata,
  m_axis_0_tready,
  m_axis_0_tvalid,
  m_axis_0_tdata
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aclk, ASSOCIATED_BUSIF m_axis_0:m_axis_1:m_axis_2:m_axis_3:m_axis_4:m_axis_5:s_axilite, ASSOCIATED_RESET aresetn, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 aclk CLK" *)
input wire aclk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME aresetn, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 aresetn RST" *)
input wire aresetn;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWREADY" *)
output wire awready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWVALID" *)
input wire awvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWADDR" *)
input wire [15 : 0] awaddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite AWPROT" *)
input wire [2 : 0] awprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WREADY" *)
output wire wready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WVALID" *)
input wire wvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WDATA" *)
input wire [31 : 0] wdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite WSTRB" *)
input wire [3 : 0] wstrb;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BREADY" *)
input wire bready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BVALID" *)
output wire bvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite BRESP" *)
output wire [1 : 0] bresp;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARREADY" *)
output wire arready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARVALID" *)
input wire arvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARADDR" *)
input wire [15 : 0] araddr;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite ARPROT" *)
input wire [2 : 0] arprot;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RREADY" *)
input wire rready;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RVALID" *)
output wire rvalid;
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RRESP" *)
output wire [1 : 0] rresp;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axilite, DATA_WIDTH 32, PROTOCOL AXI4LITE, FREQ_HZ 100000000.000000, ID_WIDTH 0, ADDR_WIDTH 16, AWUSER_WIDTH 0, ARUSER_WIDTH 0, WUSER_WIDTH 0, RUSER_WIDTH 0, BUSER_WIDTH 0, READ_WRITE_MODE READ_WRITE, HAS_BURST 0, HAS_LOCK 0, HAS_PROT 1, HAS_CACHE 0, HAS_QOS 0, HAS_REGION 0, HAS_WSTRB 1, HAS_BRESP 1, HAS_RRESP 1, SUPPORTS_NARROW_BURST 0, NUM_READ_OUTSTANDING 1, NUM_WRITE_OUTSTANDING 1, MAX_BURST_LENGTH 1, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, NUM_READ_THREADS 1, NUM_W\
RITE_THREADS 1, RUSER_BITS_PER_BYTE 0, WUSER_BITS_PER_BYTE 0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axilite RDATA" *)
output wire [31 : 0] rdata;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TREADY" *)
input wire m_axis_0_tready;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TVALID" *)
output wire m_axis_0_tvalid;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME m_axis_0, TDATA_NUM_BYTES 16, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 TDATA" *)
output wire [127 : 0] m_axis_0_tdata;

  memstream #(
    .CONFIG_EN(1'B1),
    .NSTREAMS(1),
    .MEM_DEPTH(4096),
    .MEM_WIDTH(128),
    .MEM_INIT("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/"),
    .RAM_STYLE("block"),
    .STRM0_WIDTH(128),
    .STRM1_WIDTH(32),
    .STRM2_WIDTH(32),
    .STRM3_WIDTH(32),
    .STRM4_WIDTH(32),
    .STRM5_WIDTH(32),
    .STRM0_DEPTH(4096),
    .STRM1_DEPTH(2304),
    .STRM2_DEPTH(2304),
    .STRM3_DEPTH(2304),
    .STRM4_DEPTH(2304),
    .STRM5_DEPTH(2304),
    .STRM0_OFFSET(0),
    .STRM1_OFFSET(2304),
    .STRM2_OFFSET(4608),
    .STRM3_OFFSET(6912),
    .STRM4_OFFSET(9216),
    .STRM5_OFFSET(11520),
    .AXILITE_ADDR_WIDTH(16)
  ) inst (
    .aclk(aclk),
    .aresetn(aresetn),
    .awready(awready),
    .awvalid(awvalid),
    .awaddr(awaddr),
    .awprot(awprot),
    .wready(wready),
    .wvalid(wvalid),
    .wdata(wdata),
    .wstrb(wstrb),
    .bready(bready),
    .bvalid(bvalid),
    .bresp(bresp),
    .arready(arready),
    .arvalid(arvalid),
    .araddr(araddr),
    .arprot(arprot),
    .rready(rready),
    .rvalid(rvalid),
    .rresp(rresp),
    .rdata(rdata),
    .m_axis_0_afull(1'B0),
    .m_axis_0_tready(m_axis_0_tready),
    .m_axis_0_tvalid(m_axis_0_tvalid),
    .m_axis_0_tdata(m_axis_0_tdata),
    .m_axis_1_afull(1'B0),
    .m_axis_1_tready(1'B1),
    .m_axis_1_tvalid(),
    .m_axis_1_tdata(),
    .m_axis_2_afull(1'B0),
    .m_axis_2_tready(1'B1),
    .m_axis_2_tvalid(),
    .m_axis_2_tdata(),
    .m_axis_3_afull(1'B0),
    .m_axis_3_tready(1'B1),
    .m_axis_3_tvalid(),
    .m_axis_3_tdata(),
    .m_axis_4_afull(1'B0),
    .m_axis_4_tready(1'B1),
    .m_axis_4_tvalid(),
    .m_axis_4_tdata(),
    .m_axis_5_afull(1'B0),
    .m_axis_5_tready(1'B1),
    .m_axis_5_tvalid(),
    .m_axis_5_tdata()
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccYC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccYC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccYC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccYC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccYC_rom Thresholding_Batch_0_Thresholding_BatccYC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actocq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actocq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actocq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actocq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actocq_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actocq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_Batch.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module Thresholding_Batch_2_Thresholding_Batch (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state5 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [15:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [5:0] threshs_m_thresholds_13_address0;
reg    threshs_m_thresholds_13_ce0;
wire   [17:0] threshs_m_thresholds_13_q0;
wire   [5:0] threshs_m_thresholds_12_address0;
reg    threshs_m_thresholds_12_ce0;
wire   [17:0] threshs_m_thresholds_12_q0;
wire   [5:0] threshs_m_thresholds_7_address0;
reg    threshs_m_thresholds_7_ce0;
wire   [17:0] threshs_m_thresholds_7_q0;
wire   [5:0] threshs_m_thresholds_6_address0;
reg    threshs_m_thresholds_6_ce0;
wire   [17:0] threshs_m_thresholds_6_q0;
wire   [5:0] threshs_m_thresholds_5_address0;
reg    threshs_m_thresholds_5_ce0;
wire   [17:0] threshs_m_thresholds_5_q0;
wire   [5:0] threshs_m_thresholds_4_address0;
reg    threshs_m_thresholds_4_ce0;
wire   [17:0] threshs_m_thresholds_4_q0;
wire   [5:0] threshs_m_thresholds_3_address0;
reg    threshs_m_thresholds_3_ce0;
wire   [16:0] threshs_m_thresholds_3_q0;
wire   [5:0] threshs_m_thresholds_2_address0;
reg    threshs_m_thresholds_2_ce0;
wire   [16:0] threshs_m_thresholds_2_q0;
wire   [5:0] threshs_m_thresholds_1_address0;
reg    threshs_m_thresholds_1_ce0;
wire   [16:0] threshs_m_thresholds_1_q0;
wire   [5:0] threshs_m_thresholds_address0;
reg    threshs_m_thresholds_ce0;
wire   [16:0] threshs_m_thresholds_q0;
wire   [5:0] threshs_m_thresholds_11_address0;
reg    threshs_m_thresholds_11_ce0;
wire   [16:0] threshs_m_thresholds_11_q0;
wire   [5:0] threshs_m_thresholds_10_address0;
reg    threshs_m_thresholds_10_ce0;
wire   [16:0] threshs_m_thresholds_10_q0;
wire   [5:0] threshs_m_thresholds_9_address0;
reg    threshs_m_thresholds_9_ce0;
wire   [16:0] threshs_m_thresholds_9_q0;
wire   [5:0] threshs_m_thresholds_8_address0;
reg    threshs_m_thresholds_8_ce0;
wire   [16:0] threshs_m_thresholds_8_q0;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln221_fu_299_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter2;
reg   [0:0] icmp_ln221_reg_686;
reg   [0:0] icmp_ln221_reg_686_pp0_iter1_reg;
reg   [31:0] nf_assign_reg_277;
reg   [15:0] i_0_reg_288;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
reg    ap_block_state4_io;
reg    ap_block_pp0_stage0_11001;
wire   [15:0] i_fu_305_p2;
reg  signed [15:0] tmp_V_1_reg_695;
wire   [31:0] nf_1_fu_341_p3;
wire   [0:0] icmp_ln899_fu_355_p2;
reg   [0:0] icmp_ln899_reg_776;
wire   [0:0] icmp_ln899_1_fu_361_p2;
reg   [0:0] icmp_ln899_1_reg_781;
wire   [0:0] icmp_ln899_2_fu_367_p2;
reg   [0:0] icmp_ln899_2_reg_786;
wire   [0:0] icmp_ln899_3_fu_373_p2;
reg   [0:0] icmp_ln899_3_reg_791;
wire   [0:0] icmp_ln899_4_fu_379_p2;
reg   [0:0] icmp_ln899_4_reg_796;
wire   [0:0] icmp_ln899_5_fu_385_p2;
reg   [0:0] icmp_ln899_5_reg_801;
wire   [0:0] icmp_ln899_6_fu_391_p2;
reg   [0:0] icmp_ln899_6_reg_806;
wire   [0:0] icmp_ln899_10_fu_445_p2;
reg   [0:0] icmp_ln899_10_reg_811;
wire   [0:0] icmp_ln899_11_fu_451_p2;
reg   [0:0] icmp_ln899_11_reg_816;
wire   [0:0] icmp_ln899_12_fu_457_p2;
reg   [0:0] icmp_ln899_12_reg_821;
wire   [0:0] icmp_ln899_13_fu_463_p2;
reg   [0:0] icmp_ln899_13_reg_826;
wire   [1:0] add_ln700_7_fu_475_p2;
reg   [1:0] add_ln700_7_reg_831;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
wire   [63:0] zext_ln142_fu_311_p1;
reg    ap_block_pp0_stage0_01001;
wire   [31:0] nf_fu_329_p2;
wire   [0:0] icmp_ln235_fu_335_p2;
wire  signed [17:0] sext_ln68_fu_349_p1;
wire  signed [16:0] sext_ln137_fu_352_p1;
wire   [0:0] icmp_ln899_7_fu_397_p2;
wire   [0:0] xor_ln899_7_fu_403_p2;
wire   [0:0] icmp_ln899_8_fu_413_p2;
wire   [0:0] xor_ln899_8_fu_419_p2;
wire   [0:0] icmp_ln899_9_fu_429_p2;
wire   [0:0] xor_ln899_9_fu_435_p2;
wire   [1:0] zext_ln142_8_fu_425_p1;
wire   [1:0] zext_ln142_9_fu_441_p1;
wire   [1:0] add_ln700_6_fu_469_p2;
wire   [1:0] zext_ln142_7_fu_409_p1;
wire   [0:0] xor_ln899_fu_481_p2;
wire   [0:0] xor_ln899_1_fu_494_p2;
wire   [0:0] xor_ln899_2_fu_503_p2;
wire   [0:0] xor_ln899_3_fu_512_p2;
wire   [0:0] xor_ln899_4_fu_521_p2;
wire   [0:0] xor_ln899_5_fu_530_p2;
wire   [0:0] xor_ln899_6_fu_539_p2;
wire   [0:0] xor_ln899_10_fu_548_p2;
wire   [0:0] xor_ln899_11_fu_557_p2;
wire   [0:0] xor_ln899_12_fu_566_p2;
wire   [0:0] xor_ln899_13_fu_575_p2;
wire   [1:0] zext_ln142_1_fu_499_p1;
wire   [1:0] zext_ln142_2_fu_508_p1;
wire   [1:0] add_ln700_fu_584_p2;
wire   [3:0] zext_ln700_1_fu_590_p1;
wire   [3:0] select_ln700_fu_486_p3;
wire   [1:0] zext_ln142_3_fu_517_p1;
wire   [1:0] zext_ln142_4_fu_526_p1;
wire   [1:0] add_ln700_2_fu_600_p2;
wire   [1:0] zext_ln142_5_fu_535_p1;
wire   [1:0] zext_ln142_6_fu_544_p1;
wire   [1:0] add_ln700_3_fu_610_p2;
wire   [2:0] zext_ln700_3_fu_616_p1;
wire   [2:0] zext_ln700_2_fu_606_p1;
wire   [2:0] add_ln700_4_fu_620_p2;
wire   [3:0] zext_ln700_4_fu_626_p1;
wire   [3:0] add_ln700_1_fu_594_p2;
wire   [1:0] zext_ln142_10_fu_553_p1;
wire   [1:0] zext_ln142_11_fu_562_p1;
wire   [1:0] add_ln700_8_fu_639_p2;
wire   [1:0] zext_ln142_12_fu_571_p1;
wire   [1:0] zext_ln700_fu_580_p1;
wire   [1:0] add_ln700_9_fu_649_p2;
wire   [2:0] zext_ln700_7_fu_655_p1;
wire   [2:0] zext_ln700_6_fu_645_p1;
wire   [2:0] add_ln700_10_fu_659_p2;
wire   [2:0] zext_ln700_5_fu_636_p1;
wire   [2:0] add_ln700_11_fu_665_p2;
wire   [3:0] zext_ln700_8_fu_671_p1;
wire   [3:0] add_ln700_5_fu_630_p2;
wire   [3:0] tmp_V_fu_675_p2;
wire    ap_CS_fsm_state5;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

Thresholding_Batch_2_Thresholding_Batcbkb #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_13_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_13_address0),
    .ce0(threshs_m_thresholds_13_ce0),
    .q0(threshs_m_thresholds_13_q0)
);

Thresholding_Batch_2_Thresholding_Batccud #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_12_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_12_address0),
    .ce0(threshs_m_thresholds_12_ce0),
    .q0(threshs_m_thresholds_12_q0)
);

Thresholding_Batch_2_Thresholding_BatcdEe #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_7_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_7_address0),
    .ce0(threshs_m_thresholds_7_ce0),
    .q0(threshs_m_thresholds_7_q0)
);

Thresholding_Batch_2_Thresholding_BatceOg #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_6_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_6_address0),
    .ce0(threshs_m_thresholds_6_ce0),
    .q0(threshs_m_thresholds_6_q0)
);

Thresholding_Batch_2_Thresholding_BatcfYi #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_5_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_5_address0),
    .ce0(threshs_m_thresholds_5_ce0),
    .q0(threshs_m_thresholds_5_q0)
);

Thresholding_Batch_2_Thresholding_Batcg8j #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_4_address0),
    .ce0(threshs_m_thresholds_4_ce0),
    .q0(threshs_m_thresholds_4_q0)
);

Thresholding_Batch_2_Thresholding_Batchbi #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_3_address0),
    .ce0(threshs_m_thresholds_3_ce0),
    .q0(threshs_m_thresholds_3_q0)
);

Thresholding_Batch_2_Thresholding_Batcibs #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_2_address0),
    .ce0(threshs_m_thresholds_2_ce0),
    .q0(threshs_m_thresholds_2_q0)
);

Thresholding_Batch_2_Thresholding_BatcjbC #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_1_address0),
    .ce0(threshs_m_thresholds_1_ce0),
    .q0(threshs_m_thresholds_1_q0)
);

Thresholding_Batch_2_Thresholding_BatckbM #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_address0),
    .ce0(threshs_m_thresholds_ce0),
    .q0(threshs_m_thresholds_q0)
);

Thresholding_Batch_2_Thresholding_BatclbW #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_11_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_11_address0),
    .ce0(threshs_m_thresholds_11_ce0),
    .q0(threshs_m_thresholds_11_q0)
);

Thresholding_Batch_2_Thresholding_Batcmb6 #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_10_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_10_address0),
    .ce0(threshs_m_thresholds_10_ce0),
    .q0(threshs_m_thresholds_10_q0)
);

Thresholding_Batch_2_Thresholding_Batcncg #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_9_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_9_address0),
    .ce0(threshs_m_thresholds_9_ce0),
    .q0(threshs_m_thresholds_9_q0)
);

Thresholding_Batch_2_Thresholding_Batcocq #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_8_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_8_address0),
    .ce0(threshs_m_thresholds_8_ce0),
    .q0(threshs_m_thresholds_8_q0)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_299_p2 == 1'd0))) begin
        i_0_reg_288 <= i_fu_305_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_reg_288 <= 16'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_299_p2 == 1'd0))) begin
        nf_assign_reg_277 <= nf_1_fu_341_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        nf_assign_reg_277 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_reg_686 == 1'd0))) begin
        add_ln700_7_reg_831 <= add_ln700_7_fu_475_p2;
        icmp_ln899_10_reg_811 <= icmp_ln899_10_fu_445_p2;
        icmp_ln899_11_reg_816 <= icmp_ln899_11_fu_451_p2;
        icmp_ln899_12_reg_821 <= icmp_ln899_12_fu_457_p2;
        icmp_ln899_13_reg_826 <= icmp_ln899_13_fu_463_p2;
        icmp_ln899_1_reg_781 <= icmp_ln899_1_fu_361_p2;
        icmp_ln899_2_reg_786 <= icmp_ln899_2_fu_367_p2;
        icmp_ln899_3_reg_791 <= icmp_ln899_3_fu_373_p2;
        icmp_ln899_4_reg_796 <= icmp_ln899_4_fu_379_p2;
        icmp_ln899_5_reg_801 <= icmp_ln899_5_fu_385_p2;
        icmp_ln899_6_reg_806 <= icmp_ln899_6_fu_391_p2;
        icmp_ln899_reg_776 <= icmp_ln899_fu_355_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        icmp_ln221_reg_686 <= icmp_ln221_fu_299_p2;
        icmp_ln221_reg_686_pp0_iter1_reg <= icmp_ln221_reg_686;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_299_p2 == 1'd0))) begin
        tmp_V_1_reg_695 <= in_V_V_TDATA;
    end
end

always @ (*) begin
    if ((icmp_ln221_fu_299_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state5) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state5)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln221_fu_299_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_299_p2 == 1'd0))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln221_reg_686_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_reg_686_pp0_iter1_reg == 1'd0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_10_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_10_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_11_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_11_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_12_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_12_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_13_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_13_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_1_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_1_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_2_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_2_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_3_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_3_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_4_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_4_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_5_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_5_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_6_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_6_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_7_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_7_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_8_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_8_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_9_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_9_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_299_p2 == 1'd1)) & ~((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_299_p2 == 1'd1)))) begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln700_10_fu_659_p2 = (zext_ln700_7_fu_655_p1 + zext_ln700_6_fu_645_p1);

assign add_ln700_11_fu_665_p2 = (add_ln700_10_fu_659_p2 + zext_ln700_5_fu_636_p1);

assign add_ln700_1_fu_594_p2 = (zext_ln700_1_fu_590_p1 + select_ln700_fu_486_p3);

assign add_ln700_2_fu_600_p2 = (zext_ln142_3_fu_517_p1 + zext_ln142_4_fu_526_p1);

assign add_ln700_3_fu_610_p2 = (zext_ln142_5_fu_535_p1 + zext_ln142_6_fu_544_p1);

assign add_ln700_4_fu_620_p2 = (zext_ln700_3_fu_616_p1 + zext_ln700_2_fu_606_p1);

assign add_ln700_5_fu_630_p2 = (zext_ln700_4_fu_626_p1 + add_ln700_1_fu_594_p2);

assign add_ln700_6_fu_469_p2 = (zext_ln142_8_fu_425_p1 + zext_ln142_9_fu_441_p1);

assign add_ln700_7_fu_475_p2 = (add_ln700_6_fu_469_p2 + zext_ln142_7_fu_409_p1);

assign add_ln700_8_fu_639_p2 = (zext_ln142_10_fu_553_p1 + zext_ln142_11_fu_562_p1);

assign add_ln700_9_fu_649_p2 = (zext_ln142_12_fu_571_p1 + zext_ln700_fu_580_p1);

assign add_ln700_fu_584_p2 = (zext_ln142_1_fu_499_p1 + zext_ln142_2_fu_508_p1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state5 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_299_p2 == 1'd0));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_block_state4_io)) | ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_299_p2 == 1'd0)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_block_state4_io)) | ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_299_p2 == 1'd0)));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = ((in_V_V_TVALID == 1'b0) & (icmp_ln221_fu_299_p2 == 1'd0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state4_io = ((out_V_V_TREADY == 1'b0) & (icmp_ln221_reg_686_pp0_iter1_reg == 1'd0));
end

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign i_fu_305_p2 = (i_0_reg_288 + 16'd1);

assign icmp_ln221_fu_299_p2 = ((i_0_reg_288 == 16'd50176) ? 1'b1 : 1'b0);

assign icmp_ln235_fu_335_p2 = ((nf_fu_329_p2 == 32'd64) ? 1'b1 : 1'b0);

assign icmp_ln899_10_fu_445_p2 = (($signed(sext_ln137_fu_352_p1) < $signed(threshs_m_thresholds_11_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_11_fu_451_p2 = (($signed(sext_ln137_fu_352_p1) < $signed(threshs_m_thresholds_10_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_12_fu_457_p2 = (($signed(sext_ln137_fu_352_p1) < $signed(threshs_m_thresholds_9_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_13_fu_463_p2 = (($signed(sext_ln137_fu_352_p1) < $signed(threshs_m_thresholds_8_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_1_fu_361_p2 = (($signed(sext_ln68_fu_349_p1) < $signed(threshs_m_thresholds_12_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_2_fu_367_p2 = (($signed(sext_ln68_fu_349_p1) < $signed(threshs_m_thresholds_7_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_3_fu_373_p2 = (($signed(sext_ln68_fu_349_p1) < $signed(threshs_m_thresholds_6_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_4_fu_379_p2 = (($signed(sext_ln68_fu_349_p1) < $signed(threshs_m_thresholds_5_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_5_fu_385_p2 = (($signed(sext_ln68_fu_349_p1) < $signed(threshs_m_thresholds_4_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_6_fu_391_p2 = (($signed(sext_ln137_fu_352_p1) < $signed(threshs_m_thresholds_3_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_7_fu_397_p2 = (($signed(sext_ln137_fu_352_p1) < $signed(threshs_m_thresholds_2_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_8_fu_413_p2 = (($signed(sext_ln137_fu_352_p1) < $signed(threshs_m_thresholds_1_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_9_fu_429_p2 = (($signed(sext_ln137_fu_352_p1) < $signed(threshs_m_thresholds_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_fu_355_p2 = (($signed(sext_ln68_fu_349_p1) < $signed(threshs_m_thresholds_13_q0)) ? 1'b1 : 1'b0);

assign nf_1_fu_341_p3 = ((icmp_ln235_fu_335_p2[0:0] === 1'b1) ? 32'd0 : nf_fu_329_p2);

assign nf_fu_329_p2 = (nf_assign_reg_277 + 32'd1);

assign out_V_V_TDATA = tmp_V_fu_675_p2;

assign select_ln700_fu_486_p3 = ((xor_ln899_fu_481_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign sext_ln137_fu_352_p1 = tmp_V_1_reg_695;

assign sext_ln68_fu_349_p1 = tmp_V_1_reg_695;

assign threshs_m_thresholds_10_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_11_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_12_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_13_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_1_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_2_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_3_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_4_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_5_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_6_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_7_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_8_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_9_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_address0 = zext_ln142_fu_311_p1;

assign tmp_V_fu_675_p2 = (zext_ln700_8_fu_671_p1 + add_ln700_5_fu_630_p2);

assign xor_ln899_10_fu_548_p2 = (icmp_ln899_10_reg_811 ^ 1'd1);

assign xor_ln899_11_fu_557_p2 = (icmp_ln899_11_reg_816 ^ 1'd1);

assign xor_ln899_12_fu_566_p2 = (icmp_ln899_12_reg_821 ^ 1'd1);

assign xor_ln899_13_fu_575_p2 = (icmp_ln899_13_reg_826 ^ 1'd1);

assign xor_ln899_1_fu_494_p2 = (icmp_ln899_1_reg_781 ^ 1'd1);

assign xor_ln899_2_fu_503_p2 = (icmp_ln899_2_reg_786 ^ 1'd1);

assign xor_ln899_3_fu_512_p2 = (icmp_ln899_3_reg_791 ^ 1'd1);

assign xor_ln899_4_fu_521_p2 = (icmp_ln899_4_reg_796 ^ 1'd1);

assign xor_ln899_5_fu_530_p2 = (icmp_ln899_5_reg_801 ^ 1'd1);

assign xor_ln899_6_fu_539_p2 = (icmp_ln899_6_reg_806 ^ 1'd1);

assign xor_ln899_7_fu_403_p2 = (icmp_ln899_7_fu_397_p2 ^ 1'd1);

assign xor_ln899_8_fu_419_p2 = (icmp_ln899_8_fu_413_p2 ^ 1'd1);

assign xor_ln899_9_fu_435_p2 = (icmp_ln899_9_fu_429_p2 ^ 1'd1);

assign xor_ln899_fu_481_p2 = (icmp_ln899_reg_776 ^ 1'd1);

assign zext_ln142_10_fu_553_p1 = xor_ln899_10_fu_548_p2;

assign zext_ln142_11_fu_562_p1 = xor_ln899_11_fu_557_p2;

assign zext_ln142_12_fu_571_p1 = xor_ln899_12_fu_566_p2;

assign zext_ln142_1_fu_499_p1 = xor_ln899_1_fu_494_p2;

assign zext_ln142_2_fu_508_p1 = xor_ln899_2_fu_503_p2;

assign zext_ln142_3_fu_517_p1 = xor_ln899_3_fu_512_p2;

assign zext_ln142_4_fu_526_p1 = xor_ln899_4_fu_521_p2;

assign zext_ln142_5_fu_535_p1 = xor_ln899_5_fu_530_p2;

assign zext_ln142_6_fu_544_p1 = xor_ln899_6_fu_539_p2;

assign zext_ln142_7_fu_409_p1 = xor_ln899_7_fu_403_p2;

assign zext_ln142_8_fu_425_p1 = xor_ln899_8_fu_419_p2;

assign zext_ln142_9_fu_441_p1 = xor_ln899_9_fu_435_p2;

assign zext_ln142_fu_311_p1 = nf_assign_reg_277;

assign zext_ln700_1_fu_590_p1 = add_ln700_fu_584_p2;

assign zext_ln700_2_fu_606_p1 = add_ln700_2_fu_600_p2;

assign zext_ln700_3_fu_616_p1 = add_ln700_3_fu_610_p2;

assign zext_ln700_4_fu_626_p1 = add_ln700_4_fu_620_p2;

assign zext_ln700_5_fu_636_p1 = add_ln700_7_reg_831;

assign zext_ln700_6_fu_645_p1 = add_ln700_8_fu_639_p2;

assign zext_ln700_7_fu_655_p1 = add_ln700_9_fu_649_p2;

assign zext_ln700_8_fu_671_p1 = add_ln700_11_fu_665_p2;

assign zext_ln700_fu_580_p1 = xor_ln899_13_fu_575_p2;

endmodule //Thresholding_Batch_2_Thresholding_Batch
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actyd2.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actyd2_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actyd2_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actyd2(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actyd2_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actyd2_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActUhA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActUhA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActUhA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActUhA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActUhA_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActUhA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Acthbi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Acthbi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Acthbi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Acthbi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Acthbi_rom StreamingFCLayer_Batch_4_Matrix_Vector_Acthbi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcShg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcShg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcShg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcShg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcShg_rom Thresholding_Batch_0_Thresholding_BatcShg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActCeG.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActCeG_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActCeG_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActCeG(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActCeG_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActCeG_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/466a/hdl/verilog/StreamingDataWidthConverter_Batch_1_StreamingDataWidthCo_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingDataWidthConverter_Batch_1_StreamingDataWidthCo_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state4 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [95:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [23:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln370_fu_104_p2;
wire   [0:0] icmp_ln373_fu_116_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter1;
reg   [0:0] icmp_ln370_reg_162;
reg   [71:0] p_025_0_reg_61;
reg   [31:0] o_0_reg_73;
reg   [13:0] t_0_reg_84;
reg    ap_predicate_op16_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
reg    ap_block_state3_io;
reg    ap_block_pp0_stage0_11001;
wire   [13:0] t_fu_110_p2;
reg   [0:0] icmp_ln373_reg_171;
wire   [31:0] select_ln384_fu_134_p3;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg   [95:0] ap_phi_mux_p_Val2_s_phi_fu_98_p4;
wire   [95:0] ap_phi_reg_pp0_iter0_p_Val2_s_reg_95;
reg   [95:0] ap_phi_reg_pp0_iter1_p_Val2_s_reg_95;
wire   [95:0] zext_ln370_fu_142_p1;
reg    ap_block_pp0_stage0_01001;
wire   [31:0] o_fu_122_p2;
wire   [0:0] icmp_ln384_fu_128_p2;
wire    ap_CS_fsm_state4;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_86;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_condition_86)) begin
        if (((icmp_ln373_fu_116_p2 == 1'd1) & (icmp_ln370_fu_104_p2 == 1'd0))) begin
            ap_phi_reg_pp0_iter1_p_Val2_s_reg_95 <= in_V_V_TDATA;
        end else if ((1'b1 == 1'b1)) begin
            ap_phi_reg_pp0_iter1_p_Val2_s_reg_95 <= ap_phi_reg_pp0_iter0_p_Val2_s_reg_95;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln370_fu_104_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        o_0_reg_73 <= select_ln384_fu_134_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        o_0_reg_73 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln370_reg_162 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        p_025_0_reg_61 <= {{ap_phi_mux_p_Val2_s_phi_fu_98_p4[95:24]}};
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        p_025_0_reg_61 <= 72'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln370_fu_104_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        t_0_reg_84 <= t_fu_110_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        t_0_reg_84 <= 14'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln370_reg_162 <= icmp_ln370_fu_104_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln370_fu_104_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln373_reg_171 <= icmp_ln373_fu_116_p2;
    end
end

always @ (*) begin
    if ((icmp_ln370_fu_104_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln373_reg_171 == 1'd0) & (icmp_ln370_reg_162 == 1'd0))) begin
        ap_phi_mux_p_Val2_s_phi_fu_98_p4 = zext_ln370_fu_142_p1;
    end else begin
        ap_phi_mux_p_Val2_s_phi_fu_98_p4 = ap_phi_reg_pp0_iter1_p_Val2_s_reg_95;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln373_fu_116_p2 == 1'd1) & (icmp_ln370_fu_104_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op16_read_state2 == 1'b1))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln370_reg_162 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln370_reg_162 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((icmp_ln370_fu_104_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((icmp_ln370_fu_104_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_op16_read_state2 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_op16_read_state2 == 1'b1)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_block_state3_io)) | ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_op16_read_state2 == 1'b1)));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = ((in_V_V_TVALID == 1'b0) & (ap_predicate_op16_read_state2 == 1'b1));
end

always @ (*) begin
    ap_block_state3_io = ((icmp_ln370_reg_162 == 1'd0) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_86 = ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_reg_pp0_iter0_p_Val2_s_reg_95 = 'bx;

always @ (*) begin
    ap_predicate_op16_read_state2 = ((icmp_ln373_fu_116_p2 == 1'd1) & (icmp_ln370_fu_104_p2 == 1'd0));
end

assign icmp_ln370_fu_104_p2 = ((t_0_reg_84 == 14'd12800) ? 1'b1 : 1'b0);

assign icmp_ln373_fu_116_p2 = ((o_0_reg_73 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln384_fu_128_p2 = ((o_fu_122_p2 == 32'd4) ? 1'b1 : 1'b0);

assign o_fu_122_p2 = (32'd1 + o_0_reg_73);

assign out_V_V_TDATA = ap_phi_mux_p_Val2_s_phi_fu_98_p4[23:0];

assign select_ln384_fu_134_p3 = ((icmp_ln384_fu_128_p2[0:0] === 1'b1) ? 32'd0 : o_fu_122_p2);

assign t_fu_110_p2 = (t_0_reg_84 + 14'd1);

assign zext_ln370_fu_142_p1 = p_025_0_reg_61;

endmodule //StreamingDataWidthConverter_Batch_1_StreamingDataWidthCo_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbpm.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbpm_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbpm_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbpm(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbpm_rom Thresholding_Batch_0_Thresholding_Batcbpm_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActLf8.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActLf8_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActLf8_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActLf8(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActLf8_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActLf8_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_Batcbkb_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcbkb_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_Batcbkb(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_Batcbkb_rom Thresholding_Batch_2_Thresholding_Batcbkb_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActThq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActThq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActThq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActThq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActThq_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActThq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/2c22/hdl/verilog/ConvolutionInputGenerator_2_ConvolutionInputGfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module ConvolutionInputGenerator_2_ConvolutionInputGfYi #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [23 : 0]     din0,
    input  [23 : 0]     din1,
    input  [23 : 0]     din2,
    input  [23 : 0]     din3,
    input  [1 : 0]    din4,
    output [23 : 0]   dout);

// puts internal signals
wire [1 : 0]     sel;
// level 1 signals
wire [23 : 0]         mux_1_0;
wire [23 : 0]         mux_1_1;
// level 2 signals
wire [23 : 0]         mux_2_0;

assign sel = din4;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;

// output logic
assign dout = mux_2_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Activa.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingFCLayer_Batch_4_Matrix_Vector_Activa (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY,
        weight_V_V_TDATA,
        weight_V_V_TVALID,
        weight_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state7 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [31:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;
input  [127:0] weight_V_V_TDATA;
input   weight_V_V_TVALID;
output   weight_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;
reg weight_V_V_TREADY;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [6:0] threshs_m_thresholds_55_address0;
reg    threshs_m_thresholds_55_ce0;
wire   [15:0] threshs_m_thresholds_55_q0;
wire   [6:0] threshs_m_thresholds_54_address0;
reg    threshs_m_thresholds_54_ce0;
wire   [15:0] threshs_m_thresholds_54_q0;
wire   [6:0] threshs_m_thresholds_49_address0;
reg    threshs_m_thresholds_49_ce0;
wire   [15:0] threshs_m_thresholds_49_q0;
wire   [6:0] threshs_m_thresholds_48_address0;
reg    threshs_m_thresholds_48_ce0;
wire   [15:0] threshs_m_thresholds_48_q0;
wire   [6:0] threshs_m_thresholds_47_address0;
reg    threshs_m_thresholds_47_ce0;
wire   [15:0] threshs_m_thresholds_47_q0;
wire   [6:0] threshs_m_thresholds_46_address0;
reg    threshs_m_thresholds_46_ce0;
wire   [15:0] threshs_m_thresholds_46_q0;
wire   [6:0] threshs_m_thresholds_45_address0;
reg    threshs_m_thresholds_45_ce0;
wire   [15:0] threshs_m_thresholds_45_q0;
wire   [6:0] threshs_m_thresholds_44_address0;
reg    threshs_m_thresholds_44_ce0;
wire   [15:0] threshs_m_thresholds_44_q0;
wire   [6:0] threshs_m_thresholds_43_address0;
reg    threshs_m_thresholds_43_ce0;
wire   [15:0] threshs_m_thresholds_43_q0;
wire   [6:0] threshs_m_thresholds_42_address0;
reg    threshs_m_thresholds_42_ce0;
wire   [15:0] threshs_m_thresholds_42_q0;
wire   [6:0] threshs_m_thresholds_53_address0;
reg    threshs_m_thresholds_53_ce0;
wire   [15:0] threshs_m_thresholds_53_q0;
wire   [6:0] threshs_m_thresholds_52_address0;
reg    threshs_m_thresholds_52_ce0;
wire   [15:0] threshs_m_thresholds_52_q0;
wire   [6:0] threshs_m_thresholds_51_address0;
reg    threshs_m_thresholds_51_ce0;
wire   [15:0] threshs_m_thresholds_51_q0;
wire   [6:0] threshs_m_thresholds_50_address0;
reg    threshs_m_thresholds_50_ce0;
wire   [15:0] threshs_m_thresholds_50_q0;
wire   [6:0] threshs_m_thresholds_41_address0;
reg    threshs_m_thresholds_41_ce0;
wire   [15:0] threshs_m_thresholds_41_q0;
wire   [6:0] threshs_m_thresholds_40_address0;
reg    threshs_m_thresholds_40_ce0;
wire   [15:0] threshs_m_thresholds_40_q0;
wire   [6:0] threshs_m_thresholds_35_address0;
reg    threshs_m_thresholds_35_ce0;
wire   [15:0] threshs_m_thresholds_35_q0;
wire   [6:0] threshs_m_thresholds_34_address0;
reg    threshs_m_thresholds_34_ce0;
wire   [15:0] threshs_m_thresholds_34_q0;
wire   [6:0] threshs_m_thresholds_33_address0;
reg    threshs_m_thresholds_33_ce0;
wire   [15:0] threshs_m_thresholds_33_q0;
wire   [6:0] threshs_m_thresholds_32_address0;
reg    threshs_m_thresholds_32_ce0;
wire   [15:0] threshs_m_thresholds_32_q0;
wire   [6:0] threshs_m_thresholds_31_address0;
reg    threshs_m_thresholds_31_ce0;
wire   [15:0] threshs_m_thresholds_31_q0;
wire   [6:0] threshs_m_thresholds_30_address0;
reg    threshs_m_thresholds_30_ce0;
wire   [15:0] threshs_m_thresholds_30_q0;
wire   [6:0] threshs_m_thresholds_29_address0;
reg    threshs_m_thresholds_29_ce0;
wire   [15:0] threshs_m_thresholds_29_q0;
wire   [6:0] threshs_m_thresholds_28_address0;
reg    threshs_m_thresholds_28_ce0;
wire   [15:0] threshs_m_thresholds_28_q0;
wire   [6:0] threshs_m_thresholds_39_address0;
reg    threshs_m_thresholds_39_ce0;
wire   [15:0] threshs_m_thresholds_39_q0;
wire   [6:0] threshs_m_thresholds_38_address0;
reg    threshs_m_thresholds_38_ce0;
wire   [15:0] threshs_m_thresholds_38_q0;
wire   [6:0] threshs_m_thresholds_37_address0;
reg    threshs_m_thresholds_37_ce0;
wire   [15:0] threshs_m_thresholds_37_q0;
wire   [6:0] threshs_m_thresholds_36_address0;
reg    threshs_m_thresholds_36_ce0;
wire   [15:0] threshs_m_thresholds_36_q0;
wire   [6:0] threshs_m_thresholds_27_address0;
reg    threshs_m_thresholds_27_ce0;
wire   [15:0] threshs_m_thresholds_27_q0;
wire   [6:0] threshs_m_thresholds_26_address0;
reg    threshs_m_thresholds_26_ce0;
wire   [15:0] threshs_m_thresholds_26_q0;
wire   [6:0] threshs_m_thresholds_21_address0;
reg    threshs_m_thresholds_21_ce0;
wire   [15:0] threshs_m_thresholds_21_q0;
wire   [6:0] threshs_m_thresholds_20_address0;
reg    threshs_m_thresholds_20_ce0;
wire   [15:0] threshs_m_thresholds_20_q0;
wire   [6:0] threshs_m_thresholds_19_address0;
reg    threshs_m_thresholds_19_ce0;
wire   [15:0] threshs_m_thresholds_19_q0;
wire   [6:0] threshs_m_thresholds_18_address0;
reg    threshs_m_thresholds_18_ce0;
wire   [15:0] threshs_m_thresholds_18_q0;
wire   [6:0] threshs_m_thresholds_17_address0;
reg    threshs_m_thresholds_17_ce0;
wire   [15:0] threshs_m_thresholds_17_q0;
wire   [6:0] threshs_m_thresholds_16_address0;
reg    threshs_m_thresholds_16_ce0;
wire   [15:0] threshs_m_thresholds_16_q0;
wire   [6:0] threshs_m_thresholds_15_address0;
reg    threshs_m_thresholds_15_ce0;
wire   [15:0] threshs_m_thresholds_15_q0;
wire   [6:0] threshs_m_thresholds_14_address0;
reg    threshs_m_thresholds_14_ce0;
wire   [15:0] threshs_m_thresholds_14_q0;
wire   [6:0] threshs_m_thresholds_25_address0;
reg    threshs_m_thresholds_25_ce0;
wire   [15:0] threshs_m_thresholds_25_q0;
wire   [6:0] threshs_m_thresholds_24_address0;
reg    threshs_m_thresholds_24_ce0;
wire   [15:0] threshs_m_thresholds_24_q0;
wire   [6:0] threshs_m_thresholds_23_address0;
reg    threshs_m_thresholds_23_ce0;
wire   [15:0] threshs_m_thresholds_23_q0;
wire   [6:0] threshs_m_thresholds_22_address0;
reg    threshs_m_thresholds_22_ce0;
wire   [15:0] threshs_m_thresholds_22_q0;
wire   [6:0] threshs_m_thresholds_13_address0;
reg    threshs_m_thresholds_13_ce0;
wire   [15:0] threshs_m_thresholds_13_q0;
wire   [6:0] threshs_m_thresholds_12_address0;
reg    threshs_m_thresholds_12_ce0;
wire   [15:0] threshs_m_thresholds_12_q0;
wire   [6:0] threshs_m_thresholds_7_address0;
reg    threshs_m_thresholds_7_ce0;
wire   [15:0] threshs_m_thresholds_7_q0;
wire   [6:0] threshs_m_thresholds_6_address0;
reg    threshs_m_thresholds_6_ce0;
wire   [15:0] threshs_m_thresholds_6_q0;
wire   [6:0] threshs_m_thresholds_5_address0;
reg    threshs_m_thresholds_5_ce0;
wire   [15:0] threshs_m_thresholds_5_q0;
wire   [6:0] threshs_m_thresholds_4_address0;
reg    threshs_m_thresholds_4_ce0;
wire   [15:0] threshs_m_thresholds_4_q0;
wire   [6:0] threshs_m_thresholds_3_address0;
reg    threshs_m_thresholds_3_ce0;
wire   [15:0] threshs_m_thresholds_3_q0;
wire   [6:0] threshs_m_thresholds_2_address0;
reg    threshs_m_thresholds_2_ce0;
wire   [15:0] threshs_m_thresholds_2_q0;
wire   [6:0] threshs_m_thresholds_1_address0;
reg    threshs_m_thresholds_1_ce0;
wire   [15:0] threshs_m_thresholds_1_q0;
wire   [6:0] threshs_m_thresholds_address0;
reg    threshs_m_thresholds_ce0;
wire   [15:0] threshs_m_thresholds_q0;
wire   [6:0] threshs_m_thresholds_11_address0;
reg    threshs_m_thresholds_11_ce0;
wire   [15:0] threshs_m_thresholds_11_q0;
wire   [6:0] threshs_m_thresholds_10_address0;
reg    threshs_m_thresholds_10_ce0;
wire   [15:0] threshs_m_thresholds_10_q0;
wire   [6:0] threshs_m_thresholds_9_address0;
reg    threshs_m_thresholds_9_ce0;
wire   [15:0] threshs_m_thresholds_9_q0;
wire   [6:0] threshs_m_thresholds_8_address0;
reg    threshs_m_thresholds_8_ce0;
wire   [15:0] threshs_m_thresholds_8_q0;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln248_fu_1615_p2;
wire   [0:0] icmp_ln252_fu_1630_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter4;
reg   [0:0] icmp_ln289_reg_5526;
reg   [0:0] icmp_ln289_reg_5526_pp0_iter3_reg;
reg    weight_V_V_TDATA_blk_n;
reg   [13:0] i_0_reg_1459;
reg    ap_predicate_op162_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
reg    ap_block_state6_io;
reg    ap_block_pp0_stage0_11001;
wire   [13:0] i_fu_1621_p2;
wire   [31:0] inElem_V_1_fu_1835_p66;
wire   [5:0] trunc_ln321_fu_1969_p1;
wire   [0:0] icmp_ln271_fu_2296_p2;
reg   [0:0] icmp_ln271_reg_5358;
reg   [0:0] icmp_ln271_reg_5358_pp0_iter1_reg;
wire   [3:0] wgt_M_instance_0_V_fu_2302_p1;
reg  signed [3:0] wgt_M_instance_0_V_reg_5366;
reg  signed [3:0] wgt_M_instance_1_V_reg_5371;
reg  signed [3:0] wgt_M_instance_2_V_reg_5376;
reg  signed [3:0] wgt_M_instance_3_V_reg_5381;
reg  signed [3:0] wgt_M_instance_4_V_reg_5386;
reg  signed [3:0] wgt_M_instance_5_V_reg_5391;
reg  signed [3:0] wgt_M_instance_6_V_reg_5396;
reg  signed [3:0] wgt_M_instance_7_V_reg_5401;
reg  signed [3:0] wgt_M_instance_0_V_1_reg_5406;
reg  signed [3:0] wgt_M_instance_1_V_1_reg_5411;
reg  signed [3:0] wgt_M_instance_2_V_1_reg_5416;
reg  signed [3:0] wgt_M_instance_3_V_1_reg_5421;
reg  signed [3:0] wgt_M_instance_4_V_1_reg_5426;
reg  signed [3:0] wgt_M_instance_5_V_1_reg_5431;
reg  signed [3:0] wgt_M_instance_6_V_1_reg_5436;
reg  signed [3:0] wgt_M_instance_7_V_1_reg_5441;
reg  signed [3:0] wgt_M_instance_0_V_2_reg_5446;
reg  signed [3:0] wgt_M_instance_1_V_2_reg_5451;
reg  signed [3:0] wgt_M_instance_2_V_2_reg_5456;
reg  signed [3:0] wgt_M_instance_3_V_2_reg_5461;
reg  signed [3:0] wgt_M_instance_4_V_2_reg_5466;
reg  signed [3:0] wgt_M_instance_5_V_2_reg_5471;
reg  signed [3:0] wgt_M_instance_6_V_2_reg_5476;
reg  signed [3:0] wgt_M_instance_7_V_2_reg_5481;
reg  signed [3:0] wgt_M_instance_0_V_3_reg_5486;
reg  signed [3:0] wgt_M_instance_1_V_3_reg_5491;
reg  signed [3:0] wgt_M_instance_2_V_3_reg_5496;
reg  signed [3:0] wgt_M_instance_3_V_3_reg_5501;
reg  signed [3:0] wgt_M_instance_4_V_3_reg_5506;
reg  signed [3:0] wgt_M_instance_5_V_3_reg_5511;
reg  signed [3:0] wgt_M_instance_6_V_3_reg_5516;
reg  signed [3:0] wgt_M_instance_7_V_3_reg_5521;
wire   [0:0] icmp_ln289_fu_2622_p2;
reg   [0:0] icmp_ln289_reg_5526_pp0_iter1_reg;
reg   [0:0] icmp_ln289_reg_5526_pp0_iter2_reg;
wire  signed [7:0] mul_ln1352_5_fu_2779_p2;
reg  signed [7:0] mul_ln1352_5_reg_5530;
wire   [8:0] add_ln700_1_fu_2839_p2;
reg   [8:0] add_ln700_1_reg_5535;
wire   [8:0] add_ln700_3_fu_2845_p2;
reg   [8:0] add_ln700_3_reg_5540;
wire   [8:0] add_ln700_5_fu_2857_p2;
reg   [8:0] add_ln700_5_reg_5545;
wire  signed [7:0] mul_ln1352_13_fu_2931_p2;
reg  signed [7:0] mul_ln1352_13_reg_5550;
wire   [8:0] add_ln700_9_fu_2963_p2;
reg   [8:0] add_ln700_9_reg_5555;
wire   [8:0] add_ln700_11_fu_2969_p2;
reg   [8:0] add_ln700_11_reg_5560;
wire   [8:0] add_ln700_13_fu_2981_p2;
reg   [8:0] add_ln700_13_reg_5565;
wire  signed [7:0] mul_ln1352_21_fu_3055_p2;
reg  signed [7:0] mul_ln1352_21_reg_5570;
wire   [8:0] add_ln700_17_fu_3087_p2;
reg   [8:0] add_ln700_17_reg_5575;
wire   [8:0] add_ln700_19_fu_3093_p2;
reg   [8:0] add_ln700_19_reg_5580;
wire   [8:0] add_ln700_21_fu_3105_p2;
reg   [8:0] add_ln700_21_reg_5585;
wire  signed [7:0] mul_ln1352_29_fu_3179_p2;
reg  signed [7:0] mul_ln1352_29_reg_5590;
wire   [8:0] add_ln700_25_fu_3211_p2;
reg   [8:0] add_ln700_25_reg_5595;
wire   [8:0] add_ln700_27_fu_3217_p2;
reg   [8:0] add_ln700_27_reg_5600;
wire   [8:0] add_ln700_29_fu_3229_p2;
reg   [8:0] add_ln700_29_reg_5605;
wire   [0:0] icmp_ln899_fu_3543_p2;
reg   [0:0] icmp_ln899_reg_5890;
reg   [0:0] icmp_ln899_reg_5890_pp0_iter3_reg;
wire   [0:0] icmp_ln899_1_fu_3549_p2;
reg   [0:0] icmp_ln899_1_reg_5895;
reg   [0:0] icmp_ln899_1_reg_5895_pp0_iter3_reg;
wire   [0:0] icmp_ln899_2_fu_3555_p2;
reg   [0:0] icmp_ln899_2_reg_5900;
reg   [0:0] icmp_ln899_2_reg_5900_pp0_iter3_reg;
wire   [0:0] icmp_ln899_3_fu_3561_p2;
reg   [0:0] icmp_ln899_3_reg_5905;
wire   [0:0] icmp_ln899_4_fu_3567_p2;
reg   [0:0] icmp_ln899_4_reg_5910;
wire   [0:0] icmp_ln899_5_fu_3573_p2;
reg   [0:0] icmp_ln899_5_reg_5915;
wire   [0:0] icmp_ln899_6_fu_3579_p2;
reg   [0:0] icmp_ln899_6_reg_5920;
wire   [0:0] icmp_ln899_7_fu_3585_p2;
reg   [0:0] icmp_ln899_7_reg_5925;
wire   [0:0] icmp_ln899_8_fu_3591_p2;
reg   [0:0] icmp_ln899_8_reg_5930;
wire   [0:0] icmp_ln899_9_fu_3597_p2;
reg   [0:0] icmp_ln899_9_reg_5935;
wire   [0:0] icmp_ln899_10_fu_3603_p2;
reg   [0:0] icmp_ln899_10_reg_5940;
wire   [0:0] icmp_ln899_11_fu_3609_p2;
reg   [0:0] icmp_ln899_11_reg_5945;
wire   [0:0] icmp_ln899_12_fu_3615_p2;
reg   [0:0] icmp_ln899_12_reg_5950;
wire   [0:0] icmp_ln899_13_fu_3621_p2;
reg   [0:0] icmp_ln899_13_reg_5955;
wire   [0:0] icmp_ln899_14_fu_3627_p2;
reg   [0:0] icmp_ln899_14_reg_5960;
reg   [0:0] icmp_ln899_14_reg_5960_pp0_iter3_reg;
wire   [0:0] icmp_ln899_15_fu_3633_p2;
reg   [0:0] icmp_ln899_15_reg_5965;
reg   [0:0] icmp_ln899_15_reg_5965_pp0_iter3_reg;
wire   [0:0] icmp_ln899_16_fu_3639_p2;
reg   [0:0] icmp_ln899_16_reg_5970;
reg   [0:0] icmp_ln899_16_reg_5970_pp0_iter3_reg;
wire   [0:0] icmp_ln899_17_fu_3645_p2;
reg   [0:0] icmp_ln899_17_reg_5975;
wire   [0:0] icmp_ln899_18_fu_3651_p2;
reg   [0:0] icmp_ln899_18_reg_5980;
wire   [0:0] icmp_ln899_19_fu_3657_p2;
reg   [0:0] icmp_ln899_19_reg_5985;
wire   [0:0] icmp_ln899_20_fu_3663_p2;
reg   [0:0] icmp_ln899_20_reg_5990;
wire   [0:0] icmp_ln899_21_fu_3669_p2;
reg   [0:0] icmp_ln899_21_reg_5995;
wire   [0:0] icmp_ln899_22_fu_3675_p2;
reg   [0:0] icmp_ln899_22_reg_6000;
wire   [0:0] icmp_ln899_23_fu_3681_p2;
reg   [0:0] icmp_ln899_23_reg_6005;
wire   [0:0] icmp_ln899_24_fu_3687_p2;
reg   [0:0] icmp_ln899_24_reg_6010;
wire   [0:0] icmp_ln899_25_fu_3693_p2;
reg   [0:0] icmp_ln899_25_reg_6015;
wire   [0:0] icmp_ln899_26_fu_3699_p2;
reg   [0:0] icmp_ln899_26_reg_6020;
wire   [0:0] icmp_ln899_27_fu_3705_p2;
reg   [0:0] icmp_ln899_27_reg_6025;
wire   [0:0] icmp_ln899_28_fu_3711_p2;
reg   [0:0] icmp_ln899_28_reg_6030;
reg   [0:0] icmp_ln899_28_reg_6030_pp0_iter3_reg;
wire   [0:0] icmp_ln899_29_fu_3717_p2;
reg   [0:0] icmp_ln899_29_reg_6035;
reg   [0:0] icmp_ln899_29_reg_6035_pp0_iter3_reg;
wire   [0:0] icmp_ln899_30_fu_3723_p2;
reg   [0:0] icmp_ln899_30_reg_6040;
reg   [0:0] icmp_ln899_30_reg_6040_pp0_iter3_reg;
wire   [0:0] icmp_ln899_31_fu_3729_p2;
reg   [0:0] icmp_ln899_31_reg_6045;
wire   [0:0] icmp_ln899_32_fu_3735_p2;
reg   [0:0] icmp_ln899_32_reg_6050;
wire   [0:0] icmp_ln899_33_fu_3741_p2;
reg   [0:0] icmp_ln899_33_reg_6055;
wire   [0:0] icmp_ln899_34_fu_3747_p2;
reg   [0:0] icmp_ln899_34_reg_6060;
wire   [0:0] icmp_ln899_35_fu_3753_p2;
reg   [0:0] icmp_ln899_35_reg_6065;
wire   [0:0] icmp_ln899_36_fu_3759_p2;
reg   [0:0] icmp_ln899_36_reg_6070;
wire   [0:0] icmp_ln899_37_fu_3765_p2;
reg   [0:0] icmp_ln899_37_reg_6075;
wire   [0:0] icmp_ln899_38_fu_3771_p2;
reg   [0:0] icmp_ln899_38_reg_6080;
wire   [0:0] icmp_ln899_39_fu_3777_p2;
reg   [0:0] icmp_ln899_39_reg_6085;
wire   [0:0] icmp_ln899_40_fu_3783_p2;
reg   [0:0] icmp_ln899_40_reg_6090;
wire   [0:0] icmp_ln899_41_fu_3789_p2;
reg   [0:0] icmp_ln899_41_reg_6095;
wire   [0:0] icmp_ln899_42_fu_3795_p2;
reg   [0:0] icmp_ln899_42_reg_6100;
reg   [0:0] icmp_ln899_42_reg_6100_pp0_iter3_reg;
wire   [0:0] icmp_ln899_43_fu_3801_p2;
reg   [0:0] icmp_ln899_43_reg_6105;
reg   [0:0] icmp_ln899_43_reg_6105_pp0_iter3_reg;
wire   [0:0] icmp_ln899_44_fu_3807_p2;
reg   [0:0] icmp_ln899_44_reg_6110;
reg   [0:0] icmp_ln899_44_reg_6110_pp0_iter3_reg;
wire   [0:0] icmp_ln899_45_fu_3813_p2;
reg   [0:0] icmp_ln899_45_reg_6115;
wire   [0:0] icmp_ln899_46_fu_3819_p2;
reg   [0:0] icmp_ln899_46_reg_6120;
wire   [0:0] icmp_ln899_47_fu_3825_p2;
reg   [0:0] icmp_ln899_47_reg_6125;
wire   [0:0] icmp_ln899_48_fu_3831_p2;
reg   [0:0] icmp_ln899_48_reg_6130;
wire   [0:0] icmp_ln899_49_fu_3837_p2;
reg   [0:0] icmp_ln899_49_reg_6135;
wire   [0:0] icmp_ln899_50_fu_3843_p2;
reg   [0:0] icmp_ln899_50_reg_6140;
wire   [0:0] icmp_ln899_51_fu_3849_p2;
reg   [0:0] icmp_ln899_51_reg_6145;
wire   [0:0] icmp_ln899_52_fu_3855_p2;
reg   [0:0] icmp_ln899_52_reg_6150;
wire   [0:0] icmp_ln899_53_fu_3861_p2;
reg   [0:0] icmp_ln899_53_reg_6155;
wire   [0:0] icmp_ln899_54_fu_3867_p2;
reg   [0:0] icmp_ln899_54_reg_6160;
wire   [0:0] icmp_ln899_55_fu_3873_p2;
reg   [0:0] icmp_ln899_55_reg_6165;
wire   [2:0] add_ln700_36_fu_3998_p2;
reg   [2:0] add_ln700_36_reg_6170;
wire   [2:0] add_ln700_43_fu_4046_p2;
reg   [2:0] add_ln700_43_reg_6175;
wire   [2:0] add_ln700_49_fu_4171_p2;
reg   [2:0] add_ln700_49_reg_6180;
wire   [2:0] add_ln700_56_fu_4219_p2;
reg   [2:0] add_ln700_56_reg_6185;
wire   [2:0] add_ln700_62_fu_4344_p2;
reg   [2:0] add_ln700_62_reg_6190;
wire   [2:0] add_ln700_69_fu_4392_p2;
reg   [2:0] add_ln700_69_reg_6195;
wire   [2:0] add_ln700_75_fu_4517_p2;
reg   [2:0] add_ln700_75_reg_6200;
wire   [2:0] add_ln700_82_fu_4565_p2;
reg   [2:0] add_ln700_82_reg_6205;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
wire   [31:0] ap_phi_reg_pp0_iter0_act_m_val_V_reg_1470;
reg   [31:0] ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470;
wire   [63:0] zext_ln142_fu_3238_p1;
reg   [15:0] accu_V_0_0_0_fu_432;
wire   [15:0] accu_0_0_V_fu_3397_p2;
reg   [15:0] accu_V_0_1_0_fu_436;
wire   [15:0] accu_0_1_V_fu_3437_p2;
reg   [15:0] accu_V_0_2_0_fu_440;
wire   [15:0] accu_0_2_V_fu_3477_p2;
reg   [15:0] accu_V_0_3_0_fu_444;
wire   [15:0] accu_0_3_V_fu_3517_p2;
reg   [31:0] sf_1_fu_448;
wire   [31:0] sf_fu_2616_p2;
reg   [31:0] tmp_V_fu_452;
reg   [31:0] tmp_V_1_fu_456;
reg   [31:0] tmp_V_2_fu_460;
reg   [31:0] tmp_V_4_fu_464;
reg   [31:0] tmp_V_5_fu_468;
reg   [31:0] tmp_V_6_fu_472;
reg   [31:0] tmp_V_7_fu_476;
reg   [31:0] tmp_V_8_fu_480;
reg   [31:0] tmp_V_9_fu_484;
reg   [31:0] tmp_V_10_fu_488;
reg   [31:0] tmp_V_11_fu_492;
reg   [31:0] tmp_V_12_fu_496;
reg   [31:0] tmp_V_13_fu_500;
reg   [31:0] tmp_V_14_fu_504;
reg   [31:0] tmp_V_15_fu_508;
reg   [31:0] tmp_V_16_fu_512;
reg   [31:0] tmp_V_17_fu_516;
reg   [31:0] tmp_V_18_fu_520;
reg   [31:0] tmp_V_19_fu_524;
reg   [31:0] tmp_V_20_fu_528;
reg   [31:0] tmp_V_21_fu_532;
reg   [31:0] tmp_V_22_fu_536;
reg   [31:0] tmp_V_23_fu_540;
reg   [31:0] tmp_V_24_fu_544;
reg   [31:0] tmp_V_25_fu_548;
reg   [31:0] tmp_V_26_fu_552;
reg   [31:0] tmp_V_27_fu_556;
reg   [31:0] tmp_V_28_fu_560;
reg   [31:0] tmp_V_29_fu_564;
reg   [31:0] tmp_V_30_fu_568;
reg   [31:0] tmp_V_31_fu_572;
reg   [31:0] tmp_V_32_fu_576;
reg   [31:0] tmp_V_33_fu_580;
reg   [31:0] tmp_V_34_fu_584;
reg   [31:0] tmp_V_35_fu_588;
reg   [31:0] tmp_V_36_fu_592;
reg   [31:0] tmp_V_37_fu_596;
reg   [31:0] tmp_V_38_fu_600;
reg   [31:0] tmp_V_39_fu_604;
reg   [31:0] tmp_V_40_fu_608;
reg   [31:0] tmp_V_41_fu_612;
reg   [31:0] tmp_V_42_fu_616;
reg   [31:0] tmp_V_43_fu_620;
reg   [31:0] tmp_V_44_fu_624;
reg   [31:0] tmp_V_45_fu_628;
reg   [31:0] tmp_V_46_fu_632;
reg   [31:0] tmp_V_47_fu_636;
reg   [31:0] tmp_V_48_fu_640;
reg   [31:0] tmp_V_49_fu_644;
reg   [31:0] tmp_V_50_fu_648;
reg   [31:0] tmp_V_51_fu_652;
reg   [31:0] tmp_V_52_fu_656;
reg   [31:0] tmp_V_53_fu_660;
reg   [31:0] tmp_V_54_fu_664;
reg   [31:0] tmp_V_55_fu_668;
reg   [31:0] tmp_V_56_fu_672;
reg   [31:0] tmp_V_57_fu_676;
reg   [31:0] tmp_V_58_fu_680;
reg   [31:0] tmp_V_59_fu_684;
reg   [31:0] tmp_V_60_fu_688;
reg   [31:0] tmp_V_61_fu_692;
reg   [31:0] tmp_V_62_fu_696;
reg   [31:0] tmp_V_63_fu_700;
reg   [31:0] tmp_V_64_fu_704;
reg   [31:0] nf_assign_fu_708;
wire   [31:0] select_ln301_fu_3310_p3;
reg   [31:0] ap_sig_allocacmp_nf_assign_load_1;
reg    ap_block_pp0_stage0_01001;
wire   [5:0] inElem_V_1_fu_1835_p65;
wire   [3:0] trunc_ln647_fu_2633_p1;
wire  signed [3:0] mul_ln1352_fu_2644_p0;
wire  signed [7:0] sext_ln215_1_fu_2640_p1;
wire  signed [7:0] mul_ln1352_fu_2644_p2;
wire   [3:0] arg_V_read_assign_1_fu_2654_p4;
wire  signed [3:0] mul_ln1352_1_fu_2671_p0;
wire  signed [7:0] sext_ln215_3_fu_2667_p1;
wire  signed [7:0] mul_ln1352_1_fu_2671_p2;
wire   [3:0] arg_V_read_assign_2_fu_2681_p4;
wire  signed [3:0] mul_ln1352_2_fu_2698_p0;
wire  signed [7:0] sext_ln215_5_fu_2694_p1;
wire  signed [7:0] mul_ln1352_2_fu_2698_p2;
wire   [3:0] arg_V_read_assign_3_fu_2708_p4;
wire  signed [3:0] mul_ln1352_3_fu_2725_p0;
wire  signed [7:0] sext_ln215_7_fu_2721_p1;
wire  signed [7:0] mul_ln1352_3_fu_2725_p2;
wire   [3:0] arg_V_read_assign_4_fu_2735_p4;
wire  signed [3:0] mul_ln1352_4_fu_2752_p0;
wire  signed [7:0] sext_ln215_9_fu_2748_p1;
wire  signed [7:0] mul_ln1352_4_fu_2752_p2;
wire   [3:0] arg_V_read_assign_5_fu_2762_p4;
wire  signed [3:0] mul_ln1352_5_fu_2779_p0;
wire  signed [7:0] sext_ln215_11_fu_2775_p1;
wire   [3:0] arg_V_read_assign_6_fu_2785_p4;
wire  signed [3:0] mul_ln1352_6_fu_2802_p0;
wire  signed [7:0] sext_ln215_13_fu_2798_p1;
wire  signed [7:0] mul_ln1352_6_fu_2802_p2;
wire   [3:0] arg_V_read_assign_7_fu_2812_p4;
wire  signed [3:0] mul_ln1352_7_fu_2829_p0;
wire  signed [7:0] sext_ln215_15_fu_2825_p1;
wire  signed [7:0] mul_ln1352_7_fu_2829_p2;
wire  signed [8:0] sext_ln170_4_fu_2758_p1;
wire  signed [8:0] sext_ln170_5_fu_2808_p1;
wire  signed [8:0] sext_ln170_fu_2650_p1;
wire  signed [8:0] sext_ln170_3_fu_2731_p1;
wire  signed [8:0] sext_ln700_1_fu_2835_p1;
wire  signed [8:0] sext_ln170_1_fu_2677_p1;
wire  signed [8:0] sext_ln170_2_fu_2704_p1;
wire   [8:0] add_ln700_4_fu_2851_p2;
wire  signed [3:0] mul_ln1352_8_fu_2866_p0;
wire  signed [7:0] mul_ln1352_8_fu_2866_p2;
wire  signed [3:0] mul_ln1352_9_fu_2879_p0;
wire  signed [7:0] mul_ln1352_9_fu_2879_p2;
wire  signed [3:0] mul_ln1352_10_fu_2892_p0;
wire  signed [7:0] mul_ln1352_10_fu_2892_p2;
wire  signed [3:0] mul_ln1352_11_fu_2905_p0;
wire  signed [7:0] mul_ln1352_11_fu_2905_p2;
wire  signed [3:0] mul_ln1352_12_fu_2918_p0;
wire  signed [7:0] mul_ln1352_12_fu_2918_p2;
wire  signed [3:0] mul_ln1352_13_fu_2931_p0;
wire  signed [3:0] mul_ln1352_14_fu_2940_p0;
wire  signed [7:0] mul_ln1352_14_fu_2940_p2;
wire  signed [3:0] mul_ln1352_15_fu_2953_p0;
wire  signed [7:0] mul_ln1352_15_fu_2953_p2;
wire  signed [8:0] sext_ln170_10_fu_2924_p1;
wire  signed [8:0] sext_ln170_11_fu_2946_p1;
wire  signed [8:0] sext_ln170_6_fu_2872_p1;
wire  signed [8:0] sext_ln170_9_fu_2911_p1;
wire  signed [8:0] sext_ln700_7_fu_2959_p1;
wire  signed [8:0] sext_ln170_7_fu_2885_p1;
wire  signed [8:0] sext_ln170_8_fu_2898_p1;
wire   [8:0] add_ln700_12_fu_2975_p2;
wire  signed [3:0] mul_ln1352_16_fu_2990_p0;
wire  signed [7:0] mul_ln1352_16_fu_2990_p2;
wire  signed [3:0] mul_ln1352_17_fu_3003_p0;
wire  signed [7:0] mul_ln1352_17_fu_3003_p2;
wire  signed [3:0] mul_ln1352_18_fu_3016_p0;
wire  signed [7:0] mul_ln1352_18_fu_3016_p2;
wire  signed [3:0] mul_ln1352_19_fu_3029_p0;
wire  signed [7:0] mul_ln1352_19_fu_3029_p2;
wire  signed [3:0] mul_ln1352_20_fu_3042_p0;
wire  signed [7:0] mul_ln1352_20_fu_3042_p2;
wire  signed [3:0] mul_ln1352_21_fu_3055_p0;
wire  signed [3:0] mul_ln1352_22_fu_3064_p0;
wire  signed [7:0] mul_ln1352_22_fu_3064_p2;
wire  signed [3:0] mul_ln1352_23_fu_3077_p0;
wire  signed [7:0] mul_ln1352_23_fu_3077_p2;
wire  signed [8:0] sext_ln170_16_fu_3048_p1;
wire  signed [8:0] sext_ln170_17_fu_3070_p1;
wire  signed [8:0] sext_ln170_12_fu_2996_p1;
wire  signed [8:0] sext_ln170_15_fu_3035_p1;
wire  signed [8:0] sext_ln700_13_fu_3083_p1;
wire  signed [8:0] sext_ln170_13_fu_3009_p1;
wire  signed [8:0] sext_ln170_14_fu_3022_p1;
wire   [8:0] add_ln700_20_fu_3099_p2;
wire  signed [3:0] mul_ln1352_24_fu_3114_p0;
wire  signed [7:0] mul_ln1352_24_fu_3114_p2;
wire  signed [3:0] mul_ln1352_25_fu_3127_p0;
wire  signed [7:0] mul_ln1352_25_fu_3127_p2;
wire  signed [3:0] mul_ln1352_26_fu_3140_p0;
wire  signed [7:0] mul_ln1352_26_fu_3140_p2;
wire  signed [3:0] mul_ln1352_27_fu_3153_p0;
wire  signed [7:0] mul_ln1352_27_fu_3153_p2;
wire  signed [3:0] mul_ln1352_28_fu_3166_p0;
wire  signed [7:0] mul_ln1352_28_fu_3166_p2;
wire  signed [3:0] mul_ln1352_29_fu_3179_p0;
wire  signed [3:0] mul_ln1352_30_fu_3188_p0;
wire  signed [7:0] mul_ln1352_30_fu_3188_p2;
wire  signed [3:0] mul_ln1352_31_fu_3201_p0;
wire  signed [7:0] mul_ln1352_31_fu_3201_p2;
wire  signed [8:0] sext_ln170_22_fu_3172_p1;
wire  signed [8:0] sext_ln170_23_fu_3194_p1;
wire  signed [8:0] sext_ln170_18_fu_3120_p1;
wire  signed [8:0] sext_ln170_21_fu_3159_p1;
wire  signed [8:0] sext_ln700_19_fu_3207_p1;
wire  signed [8:0] sext_ln170_19_fu_3133_p1;
wire  signed [8:0] sext_ln170_20_fu_3146_p1;
wire   [8:0] add_ln700_28_fu_3223_p2;
wire   [31:0] nf_fu_3298_p2;
wire   [0:0] icmp_ln301_fu_3304_p2;
wire  signed [15:0] sext_ln700_fu_3363_p1;
wire   [15:0] select_ln271_3_fu_3356_p3;
wire   [15:0] add_ln700_fu_3366_p2;
wire  signed [15:0] sext_ln700_2_fu_3372_p1;
wire  signed [9:0] sext_ln700_3_fu_3381_p1;
wire  signed [9:0] sext_ln700_4_fu_3384_p1;
wire   [9:0] add_ln700_6_fu_3387_p2;
wire   [15:0] add_ln700_2_fu_3375_p2;
wire  signed [15:0] sext_ln700_5_fu_3393_p1;
wire  signed [15:0] sext_ln700_6_fu_3403_p1;
wire   [15:0] select_ln271_2_fu_3349_p3;
wire   [15:0] add_ln700_8_fu_3406_p2;
wire  signed [15:0] sext_ln700_8_fu_3412_p1;
wire  signed [9:0] sext_ln700_9_fu_3421_p1;
wire  signed [9:0] sext_ln700_10_fu_3424_p1;
wire   [9:0] add_ln700_14_fu_3427_p2;
wire   [15:0] add_ln700_10_fu_3415_p2;
wire  signed [15:0] sext_ln700_11_fu_3433_p1;
wire  signed [15:0] sext_ln700_12_fu_3443_p1;
wire   [15:0] select_ln271_1_fu_3342_p3;
wire   [15:0] add_ln700_16_fu_3446_p2;
wire  signed [15:0] sext_ln700_14_fu_3452_p1;
wire  signed [9:0] sext_ln700_15_fu_3461_p1;
wire  signed [9:0] sext_ln700_16_fu_3464_p1;
wire   [9:0] add_ln700_22_fu_3467_p2;
wire   [15:0] add_ln700_18_fu_3455_p2;
wire  signed [15:0] sext_ln700_17_fu_3473_p1;
wire  signed [15:0] sext_ln700_18_fu_3483_p1;
wire   [15:0] select_ln271_fu_3335_p3;
wire   [15:0] add_ln700_24_fu_3486_p2;
wire  signed [15:0] sext_ln700_20_fu_3492_p1;
wire  signed [9:0] sext_ln700_21_fu_3501_p1;
wire  signed [9:0] sext_ln700_22_fu_3504_p1;
wire   [9:0] add_ln700_30_fu_3507_p2;
wire   [15:0] add_ln700_26_fu_3495_p2;
wire  signed [15:0] sext_ln700_23_fu_3513_p1;
wire   [0:0] xor_ln899_3_fu_3879_p2;
wire   [0:0] xor_ln899_4_fu_3888_p2;
wire   [0:0] xor_ln899_5_fu_3897_p2;
wire   [0:0] xor_ln899_6_fu_3906_p2;
wire   [0:0] xor_ln899_7_fu_3915_p2;
wire   [0:0] xor_ln899_8_fu_3924_p2;
wire   [0:0] xor_ln899_9_fu_3933_p2;
wire   [0:0] xor_ln899_10_fu_3942_p2;
wire   [0:0] xor_ln899_11_fu_3951_p2;
wire   [0:0] xor_ln899_12_fu_3960_p2;
wire   [0:0] xor_ln899_13_fu_3969_p2;
wire   [1:0] zext_ln142_3_fu_3884_p1;
wire   [1:0] zext_ln142_4_fu_3893_p1;
wire   [1:0] add_ln700_34_fu_3978_p2;
wire   [1:0] zext_ln142_5_fu_3902_p1;
wire   [1:0] zext_ln142_6_fu_3911_p1;
wire   [1:0] add_ln700_35_fu_3988_p2;
wire   [2:0] zext_ln700_3_fu_3994_p1;
wire   [2:0] zext_ln700_2_fu_3984_p1;
wire   [1:0] zext_ln142_8_fu_3929_p1;
wire   [1:0] zext_ln142_9_fu_3938_p1;
wire   [1:0] add_ln700_38_fu_4004_p2;
wire   [1:0] zext_ln142_7_fu_3920_p1;
wire   [1:0] add_ln700_39_fu_4010_p2;
wire   [1:0] zext_ln142_10_fu_3947_p1;
wire   [1:0] zext_ln142_11_fu_3956_p1;
wire   [1:0] add_ln700_40_fu_4020_p2;
wire   [1:0] zext_ln142_12_fu_3965_p1;
wire   [1:0] zext_ln700_fu_3974_p1;
wire   [1:0] add_ln700_41_fu_4030_p2;
wire   [2:0] zext_ln700_7_fu_4036_p1;
wire   [2:0] zext_ln700_6_fu_4026_p1;
wire   [2:0] add_ln700_42_fu_4040_p2;
wire   [2:0] zext_ln700_5_fu_4016_p1;
wire   [0:0] xor_ln899_17_fu_4052_p2;
wire   [0:0] xor_ln899_18_fu_4061_p2;
wire   [0:0] xor_ln899_19_fu_4070_p2;
wire   [0:0] xor_ln899_20_fu_4079_p2;
wire   [0:0] xor_ln899_21_fu_4088_p2;
wire   [0:0] xor_ln899_22_fu_4097_p2;
wire   [0:0] xor_ln899_23_fu_4106_p2;
wire   [0:0] xor_ln899_24_fu_4115_p2;
wire   [0:0] xor_ln899_25_fu_4124_p2;
wire   [0:0] xor_ln899_26_fu_4133_p2;
wire   [0:0] xor_ln899_27_fu_4142_p2;
wire   [1:0] zext_ln142_15_fu_4057_p1;
wire   [1:0] zext_ln142_16_fu_4066_p1;
wire   [1:0] add_ln700_47_fu_4151_p2;
wire   [1:0] zext_ln142_17_fu_4075_p1;
wire   [1:0] zext_ln142_18_fu_4084_p1;
wire   [1:0] add_ln700_48_fu_4161_p2;
wire   [2:0] zext_ln700_12_fu_4167_p1;
wire   [2:0] zext_ln700_11_fu_4157_p1;
wire   [1:0] zext_ln142_20_fu_4102_p1;
wire   [1:0] zext_ln142_21_fu_4111_p1;
wire   [1:0] add_ln700_51_fu_4177_p2;
wire   [1:0] zext_ln142_19_fu_4093_p1;
wire   [1:0] add_ln700_52_fu_4183_p2;
wire   [1:0] zext_ln142_22_fu_4120_p1;
wire   [1:0] zext_ln142_23_fu_4129_p1;
wire   [1:0] add_ln700_53_fu_4193_p2;
wire   [1:0] zext_ln142_24_fu_4138_p1;
wire   [1:0] zext_ln700_9_fu_4147_p1;
wire   [1:0] add_ln700_54_fu_4203_p2;
wire   [2:0] zext_ln700_16_fu_4209_p1;
wire   [2:0] zext_ln700_15_fu_4199_p1;
wire   [2:0] add_ln700_55_fu_4213_p2;
wire   [2:0] zext_ln700_14_fu_4189_p1;
wire   [0:0] xor_ln899_31_fu_4225_p2;
wire   [0:0] xor_ln899_32_fu_4234_p2;
wire   [0:0] xor_ln899_33_fu_4243_p2;
wire   [0:0] xor_ln899_34_fu_4252_p2;
wire   [0:0] xor_ln899_35_fu_4261_p2;
wire   [0:0] xor_ln899_36_fu_4270_p2;
wire   [0:0] xor_ln899_37_fu_4279_p2;
wire   [0:0] xor_ln899_38_fu_4288_p2;
wire   [0:0] xor_ln899_39_fu_4297_p2;
wire   [0:0] xor_ln899_40_fu_4306_p2;
wire   [0:0] xor_ln899_41_fu_4315_p2;
wire   [1:0] zext_ln142_27_fu_4230_p1;
wire   [1:0] zext_ln142_28_fu_4239_p1;
wire   [1:0] add_ln700_60_fu_4324_p2;
wire   [1:0] zext_ln142_29_fu_4248_p1;
wire   [1:0] zext_ln142_30_fu_4257_p1;
wire   [1:0] add_ln700_61_fu_4334_p2;
wire   [2:0] zext_ln700_21_fu_4340_p1;
wire   [2:0] zext_ln700_20_fu_4330_p1;
wire   [1:0] zext_ln142_32_fu_4275_p1;
wire   [1:0] zext_ln142_33_fu_4284_p1;
wire   [1:0] add_ln700_64_fu_4350_p2;
wire   [1:0] zext_ln142_31_fu_4266_p1;
wire   [1:0] add_ln700_65_fu_4356_p2;
wire   [1:0] zext_ln142_34_fu_4293_p1;
wire   [1:0] zext_ln142_35_fu_4302_p1;
wire   [1:0] add_ln700_66_fu_4366_p2;
wire   [1:0] zext_ln142_36_fu_4311_p1;
wire   [1:0] zext_ln700_18_fu_4320_p1;
wire   [1:0] add_ln700_67_fu_4376_p2;
wire   [2:0] zext_ln700_25_fu_4382_p1;
wire   [2:0] zext_ln700_24_fu_4372_p1;
wire   [2:0] add_ln700_68_fu_4386_p2;
wire   [2:0] zext_ln700_23_fu_4362_p1;
wire   [0:0] xor_ln899_45_fu_4398_p2;
wire   [0:0] xor_ln899_46_fu_4407_p2;
wire   [0:0] xor_ln899_47_fu_4416_p2;
wire   [0:0] xor_ln899_48_fu_4425_p2;
wire   [0:0] xor_ln899_49_fu_4434_p2;
wire   [0:0] xor_ln899_50_fu_4443_p2;
wire   [0:0] xor_ln899_51_fu_4452_p2;
wire   [0:0] xor_ln899_52_fu_4461_p2;
wire   [0:0] xor_ln899_53_fu_4470_p2;
wire   [0:0] xor_ln899_54_fu_4479_p2;
wire   [0:0] xor_ln899_55_fu_4488_p2;
wire   [1:0] zext_ln142_39_fu_4403_p1;
wire   [1:0] zext_ln142_40_fu_4412_p1;
wire   [1:0] add_ln700_73_fu_4497_p2;
wire   [1:0] zext_ln142_41_fu_4421_p1;
wire   [1:0] zext_ln142_42_fu_4430_p1;
wire   [1:0] add_ln700_74_fu_4507_p2;
wire   [2:0] zext_ln700_30_fu_4513_p1;
wire   [2:0] zext_ln700_29_fu_4503_p1;
wire   [1:0] zext_ln142_44_fu_4448_p1;
wire   [1:0] zext_ln142_45_fu_4457_p1;
wire   [1:0] add_ln700_77_fu_4523_p2;
wire   [1:0] zext_ln142_43_fu_4439_p1;
wire   [1:0] add_ln700_78_fu_4529_p2;
wire   [1:0] zext_ln142_46_fu_4466_p1;
wire   [1:0] zext_ln142_47_fu_4475_p1;
wire   [1:0] add_ln700_79_fu_4539_p2;
wire   [1:0] zext_ln142_48_fu_4484_p1;
wire   [1:0] zext_ln700_27_fu_4493_p1;
wire   [1:0] add_ln700_80_fu_4549_p2;
wire   [2:0] zext_ln700_34_fu_4555_p1;
wire   [2:0] zext_ln700_33_fu_4545_p1;
wire   [2:0] add_ln700_81_fu_4559_p2;
wire   [2:0] zext_ln700_32_fu_4535_p1;
wire   [0:0] xor_ln899_fu_4571_p2;
wire   [0:0] xor_ln899_1_fu_4584_p2;
wire   [0:0] xor_ln899_2_fu_4593_p2;
wire   [1:0] zext_ln142_1_fu_4589_p1;
wire   [1:0] zext_ln142_2_fu_4598_p1;
wire   [1:0] add_ln700_32_fu_4602_p2;
wire   [3:0] zext_ln700_1_fu_4608_p1;
wire   [3:0] select_ln700_fu_4576_p3;
wire   [3:0] zext_ln700_4_fu_4618_p1;
wire   [3:0] add_ln700_33_fu_4612_p2;
wire   [3:0] zext_ln700_8_fu_4627_p1;
wire   [3:0] add_ln700_37_fu_4621_p2;
wire   [0:0] xor_ln899_14_fu_4636_p2;
wire   [0:0] xor_ln899_15_fu_4649_p2;
wire   [0:0] xor_ln899_16_fu_4658_p2;
wire   [1:0] zext_ln142_13_fu_4654_p1;
wire   [1:0] zext_ln142_14_fu_4663_p1;
wire   [1:0] add_ln700_45_fu_4667_p2;
wire   [3:0] zext_ln700_10_fu_4673_p1;
wire   [3:0] select_ln700_1_fu_4641_p3;
wire   [3:0] zext_ln700_13_fu_4683_p1;
wire   [3:0] add_ln700_46_fu_4677_p2;
wire   [3:0] zext_ln700_17_fu_4692_p1;
wire   [3:0] add_ln700_50_fu_4686_p2;
wire   [0:0] xor_ln899_28_fu_4701_p2;
wire   [0:0] xor_ln899_29_fu_4714_p2;
wire   [0:0] xor_ln899_30_fu_4723_p2;
wire   [1:0] zext_ln142_25_fu_4719_p1;
wire   [1:0] zext_ln142_26_fu_4728_p1;
wire   [1:0] add_ln700_58_fu_4732_p2;
wire   [3:0] zext_ln700_19_fu_4738_p1;
wire   [3:0] select_ln700_2_fu_4706_p3;
wire   [3:0] zext_ln700_22_fu_4748_p1;
wire   [3:0] add_ln700_59_fu_4742_p2;
wire   [3:0] zext_ln700_26_fu_4757_p1;
wire   [3:0] add_ln700_63_fu_4751_p2;
wire   [0:0] xor_ln899_42_fu_4766_p2;
wire   [0:0] xor_ln899_43_fu_4779_p2;
wire   [0:0] xor_ln899_44_fu_4788_p2;
wire   [1:0] zext_ln142_37_fu_4784_p1;
wire   [1:0] zext_ln142_38_fu_4793_p1;
wire   [1:0] add_ln700_71_fu_4797_p2;
wire   [3:0] zext_ln700_28_fu_4803_p1;
wire   [3:0] select_ln700_3_fu_4771_p3;
wire   [3:0] zext_ln700_31_fu_4813_p1;
wire   [3:0] add_ln700_72_fu_4807_p2;
wire   [3:0] zext_ln700_35_fu_4822_p1;
wire   [3:0] add_ln700_76_fu_4816_p2;
wire   [3:0] add_ln700_83_fu_4825_p2;
wire   [3:0] add_ln700_70_fu_4760_p2;
wire   [3:0] add_ln700_57_fu_4695_p2;
wire   [3:0] add_ln700_44_fu_4630_p2;
wire    ap_CS_fsm_state7;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
end

StreamingFCLayer_Batch_4_Matrix_Vector_Actbkb #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_55_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_55_address0),
    .ce0(threshs_m_thresholds_55_ce0),
    .q0(threshs_m_thresholds_55_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actcud #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_54_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_54_address0),
    .ce0(threshs_m_thresholds_54_ce0),
    .q0(threshs_m_thresholds_54_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActdEe #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_49_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_49_address0),
    .ce0(threshs_m_thresholds_49_ce0),
    .q0(threshs_m_thresholds_49_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActeOg #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_48_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_48_address0),
    .ce0(threshs_m_thresholds_48_ce0),
    .q0(threshs_m_thresholds_48_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActfYi #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_47_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_47_address0),
    .ce0(threshs_m_thresholds_47_ce0),
    .q0(threshs_m_thresholds_47_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actg8j #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_46_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_46_address0),
    .ce0(threshs_m_thresholds_46_ce0),
    .q0(threshs_m_thresholds_46_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Acthbi #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_45_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_45_address0),
    .ce0(threshs_m_thresholds_45_ce0),
    .q0(threshs_m_thresholds_45_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actibs #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_44_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_44_address0),
    .ce0(threshs_m_thresholds_44_ce0),
    .q0(threshs_m_thresholds_44_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActjbC #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_43_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_43_address0),
    .ce0(threshs_m_thresholds_43_ce0),
    .q0(threshs_m_thresholds_43_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActkbM #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_42_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_42_address0),
    .ce0(threshs_m_thresholds_42_ce0),
    .q0(threshs_m_thresholds_42_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActlbW #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_53_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_53_address0),
    .ce0(threshs_m_thresholds_53_ce0),
    .q0(threshs_m_thresholds_53_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actmb6 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_52_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_52_address0),
    .ce0(threshs_m_thresholds_52_ce0),
    .q0(threshs_m_thresholds_52_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actncg #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_51_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_51_address0),
    .ce0(threshs_m_thresholds_51_ce0),
    .q0(threshs_m_thresholds_51_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actocq #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_50_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_50_address0),
    .ce0(threshs_m_thresholds_50_ce0),
    .q0(threshs_m_thresholds_50_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActpcA #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_41_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_41_address0),
    .ce0(threshs_m_thresholds_41_ce0),
    .q0(threshs_m_thresholds_41_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActqcK #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_40_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_40_address0),
    .ce0(threshs_m_thresholds_40_ce0),
    .q0(threshs_m_thresholds_40_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActrcU #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_35_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_35_address0),
    .ce0(threshs_m_thresholds_35_ce0),
    .q0(threshs_m_thresholds_35_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actsc4 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_34_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_34_address0),
    .ce0(threshs_m_thresholds_34_ce0),
    .q0(threshs_m_thresholds_34_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Acttde #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_33_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_33_address0),
    .ce0(threshs_m_thresholds_33_ce0),
    .q0(threshs_m_thresholds_33_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actudo #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_32_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_32_address0),
    .ce0(threshs_m_thresholds_32_ce0),
    .q0(threshs_m_thresholds_32_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actvdy #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_31_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_31_address0),
    .ce0(threshs_m_thresholds_31_ce0),
    .q0(threshs_m_thresholds_31_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActwdI #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_30_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_30_address0),
    .ce0(threshs_m_thresholds_30_ce0),
    .q0(threshs_m_thresholds_30_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActxdS #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_29_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_29_address0),
    .ce0(threshs_m_thresholds_29_ce0),
    .q0(threshs_m_thresholds_29_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actyd2 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_28_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_28_address0),
    .ce0(threshs_m_thresholds_28_ce0),
    .q0(threshs_m_thresholds_28_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Actzec #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_39_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_39_address0),
    .ce0(threshs_m_thresholds_39_ce0),
    .q0(threshs_m_thresholds_39_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActAem #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_38_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_38_address0),
    .ce0(threshs_m_thresholds_38_ce0),
    .q0(threshs_m_thresholds_38_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActBew #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_37_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_37_address0),
    .ce0(threshs_m_thresholds_37_ce0),
    .q0(threshs_m_thresholds_37_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActCeG #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_36_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_36_address0),
    .ce0(threshs_m_thresholds_36_ce0),
    .q0(threshs_m_thresholds_36_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActDeQ #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_27_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_27_address0),
    .ce0(threshs_m_thresholds_27_ce0),
    .q0(threshs_m_thresholds_27_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActEe0 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_26_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_26_address0),
    .ce0(threshs_m_thresholds_26_ce0),
    .q0(threshs_m_thresholds_26_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActFfa #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_21_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_21_address0),
    .ce0(threshs_m_thresholds_21_ce0),
    .q0(threshs_m_thresholds_21_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActGfk #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_20_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_20_address0),
    .ce0(threshs_m_thresholds_20_ce0),
    .q0(threshs_m_thresholds_20_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActHfu #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_19_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_19_address0),
    .ce0(threshs_m_thresholds_19_ce0),
    .q0(threshs_m_thresholds_19_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActIfE #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_18_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_18_address0),
    .ce0(threshs_m_thresholds_18_ce0),
    .q0(threshs_m_thresholds_18_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActJfO #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_17_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_17_address0),
    .ce0(threshs_m_thresholds_17_ce0),
    .q0(threshs_m_thresholds_17_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActKfY #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_16_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_16_address0),
    .ce0(threshs_m_thresholds_16_ce0),
    .q0(threshs_m_thresholds_16_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActLf8 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_15_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_15_address0),
    .ce0(threshs_m_thresholds_15_ce0),
    .q0(threshs_m_thresholds_15_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActMgi #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_14_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_14_address0),
    .ce0(threshs_m_thresholds_14_ce0),
    .q0(threshs_m_thresholds_14_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActNgs #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_25_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_25_address0),
    .ce0(threshs_m_thresholds_25_ce0),
    .q0(threshs_m_thresholds_25_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActOgC #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_24_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_24_address0),
    .ce0(threshs_m_thresholds_24_ce0),
    .q0(threshs_m_thresholds_24_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActPgM #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_23_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_23_address0),
    .ce0(threshs_m_thresholds_23_ce0),
    .q0(threshs_m_thresholds_23_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActQgW #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_22_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_22_address0),
    .ce0(threshs_m_thresholds_22_ce0),
    .q0(threshs_m_thresholds_22_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActRg6 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_13_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_13_address0),
    .ce0(threshs_m_thresholds_13_ce0),
    .q0(threshs_m_thresholds_13_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActShg #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_12_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_12_address0),
    .ce0(threshs_m_thresholds_12_ce0),
    .q0(threshs_m_thresholds_12_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActThq #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_7_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_7_address0),
    .ce0(threshs_m_thresholds_7_ce0),
    .q0(threshs_m_thresholds_7_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActUhA #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_6_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_6_address0),
    .ce0(threshs_m_thresholds_6_ce0),
    .q0(threshs_m_thresholds_6_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActVhK #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_5_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_5_address0),
    .ce0(threshs_m_thresholds_5_ce0),
    .q0(threshs_m_thresholds_5_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActWhU #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_4_address0),
    .ce0(threshs_m_thresholds_4_ce0),
    .q0(threshs_m_thresholds_4_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActXh4 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_3_address0),
    .ce0(threshs_m_thresholds_3_ce0),
    .q0(threshs_m_thresholds_3_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActYie #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_2_address0),
    .ce0(threshs_m_thresholds_2_ce0),
    .q0(threshs_m_thresholds_2_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_ActZio #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_1_address0),
    .ce0(threshs_m_thresholds_1_ce0),
    .q0(threshs_m_thresholds_1_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Act0iy #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_address0),
    .ce0(threshs_m_thresholds_ce0),
    .q0(threshs_m_thresholds_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Act1iI #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_11_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_11_address0),
    .ce0(threshs_m_thresholds_11_ce0),
    .q0(threshs_m_thresholds_11_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Act2iS #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_10_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_10_address0),
    .ce0(threshs_m_thresholds_10_ce0),
    .q0(threshs_m_thresholds_10_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Act3i2 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_9_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_9_address0),
    .ce0(threshs_m_thresholds_9_ce0),
    .q0(threshs_m_thresholds_9_q0)
);

StreamingFCLayer_Batch_4_Matrix_Vector_Act4jc #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_8_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_8_address0),
    .ce0(threshs_m_thresholds_8_ce0),
    .q0(threshs_m_thresholds_8_q0)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_5jm #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 32 ),
    .din5_WIDTH( 32 ),
    .din6_WIDTH( 32 ),
    .din7_WIDTH( 32 ),
    .din8_WIDTH( 32 ),
    .din9_WIDTH( 32 ),
    .din10_WIDTH( 32 ),
    .din11_WIDTH( 32 ),
    .din12_WIDTH( 32 ),
    .din13_WIDTH( 32 ),
    .din14_WIDTH( 32 ),
    .din15_WIDTH( 32 ),
    .din16_WIDTH( 32 ),
    .din17_WIDTH( 32 ),
    .din18_WIDTH( 32 ),
    .din19_WIDTH( 32 ),
    .din20_WIDTH( 32 ),
    .din21_WIDTH( 32 ),
    .din22_WIDTH( 32 ),
    .din23_WIDTH( 32 ),
    .din24_WIDTH( 32 ),
    .din25_WIDTH( 32 ),
    .din26_WIDTH( 32 ),
    .din27_WIDTH( 32 ),
    .din28_WIDTH( 32 ),
    .din29_WIDTH( 32 ),
    .din30_WIDTH( 32 ),
    .din31_WIDTH( 32 ),
    .din32_WIDTH( 32 ),
    .din33_WIDTH( 32 ),
    .din34_WIDTH( 32 ),
    .din35_WIDTH( 32 ),
    .din36_WIDTH( 32 ),
    .din37_WIDTH( 32 ),
    .din38_WIDTH( 32 ),
    .din39_WIDTH( 32 ),
    .din40_WIDTH( 32 ),
    .din41_WIDTH( 32 ),
    .din42_WIDTH( 32 ),
    .din43_WIDTH( 32 ),
    .din44_WIDTH( 32 ),
    .din45_WIDTH( 32 ),
    .din46_WIDTH( 32 ),
    .din47_WIDTH( 32 ),
    .din48_WIDTH( 32 ),
    .din49_WIDTH( 32 ),
    .din50_WIDTH( 32 ),
    .din51_WIDTH( 32 ),
    .din52_WIDTH( 32 ),
    .din53_WIDTH( 32 ),
    .din54_WIDTH( 32 ),
    .din55_WIDTH( 32 ),
    .din56_WIDTH( 32 ),
    .din57_WIDTH( 32 ),
    .din58_WIDTH( 32 ),
    .din59_WIDTH( 32 ),
    .din60_WIDTH( 32 ),
    .din61_WIDTH( 32 ),
    .din62_WIDTH( 32 ),
    .din63_WIDTH( 32 ),
    .din64_WIDTH( 6 ),
    .dout_WIDTH( 32 ))
StreamingFCLayer_5jm_U1(
    .din0(tmp_V_fu_452),
    .din1(tmp_V_1_fu_456),
    .din2(tmp_V_2_fu_460),
    .din3(tmp_V_4_fu_464),
    .din4(tmp_V_5_fu_468),
    .din5(tmp_V_6_fu_472),
    .din6(tmp_V_7_fu_476),
    .din7(tmp_V_8_fu_480),
    .din8(tmp_V_9_fu_484),
    .din9(tmp_V_10_fu_488),
    .din10(tmp_V_11_fu_492),
    .din11(tmp_V_12_fu_496),
    .din12(tmp_V_13_fu_500),
    .din13(tmp_V_14_fu_504),
    .din14(tmp_V_15_fu_508),
    .din15(tmp_V_16_fu_512),
    .din16(tmp_V_17_fu_516),
    .din17(tmp_V_18_fu_520),
    .din18(tmp_V_19_fu_524),
    .din19(tmp_V_20_fu_528),
    .din20(tmp_V_21_fu_532),
    .din21(tmp_V_22_fu_536),
    .din22(tmp_V_23_fu_540),
    .din23(tmp_V_24_fu_544),
    .din24(tmp_V_25_fu_548),
    .din25(tmp_V_26_fu_552),
    .din26(tmp_V_27_fu_556),
    .din27(tmp_V_28_fu_560),
    .din28(tmp_V_29_fu_564),
    .din29(tmp_V_30_fu_568),
    .din30(tmp_V_31_fu_572),
    .din31(tmp_V_32_fu_576),
    .din32(tmp_V_33_fu_580),
    .din33(tmp_V_34_fu_584),
    .din34(tmp_V_35_fu_588),
    .din35(tmp_V_36_fu_592),
    .din36(tmp_V_37_fu_596),
    .din37(tmp_V_38_fu_600),
    .din38(tmp_V_39_fu_604),
    .din39(tmp_V_40_fu_608),
    .din40(tmp_V_41_fu_612),
    .din41(tmp_V_42_fu_616),
    .din42(tmp_V_43_fu_620),
    .din43(tmp_V_44_fu_624),
    .din44(tmp_V_45_fu_628),
    .din45(tmp_V_46_fu_632),
    .din46(tmp_V_47_fu_636),
    .din47(tmp_V_48_fu_640),
    .din48(tmp_V_49_fu_644),
    .din49(tmp_V_50_fu_648),
    .din50(tmp_V_51_fu_652),
    .din51(tmp_V_52_fu_656),
    .din52(tmp_V_53_fu_660),
    .din53(tmp_V_54_fu_664),
    .din54(tmp_V_55_fu_668),
    .din55(tmp_V_56_fu_672),
    .din56(tmp_V_57_fu_676),
    .din57(tmp_V_58_fu_680),
    .din58(tmp_V_59_fu_684),
    .din59(tmp_V_60_fu_688),
    .din60(tmp_V_61_fu_692),
    .din61(tmp_V_62_fu_696),
    .din62(tmp_V_63_fu_700),
    .din63(tmp_V_64_fu_704),
    .din64(inElem_V_1_fu_1835_p65),
    .dout(inElem_V_1_fu_1835_p66)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U2(
    .din0(mul_ln1352_fu_2644_p0),
    .din1(wgt_M_instance_0_V_reg_5366),
    .dout(mul_ln1352_fu_2644_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U3(
    .din0(mul_ln1352_1_fu_2671_p0),
    .din1(wgt_M_instance_1_V_reg_5371),
    .dout(mul_ln1352_1_fu_2671_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U4(
    .din0(mul_ln1352_2_fu_2698_p0),
    .din1(wgt_M_instance_2_V_reg_5376),
    .dout(mul_ln1352_2_fu_2698_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U5(
    .din0(mul_ln1352_3_fu_2725_p0),
    .din1(wgt_M_instance_3_V_reg_5381),
    .dout(mul_ln1352_3_fu_2725_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U6(
    .din0(mul_ln1352_4_fu_2752_p0),
    .din1(wgt_M_instance_4_V_reg_5386),
    .dout(mul_ln1352_4_fu_2752_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U7(
    .din0(mul_ln1352_5_fu_2779_p0),
    .din1(wgt_M_instance_5_V_reg_5391),
    .dout(mul_ln1352_5_fu_2779_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U8(
    .din0(mul_ln1352_6_fu_2802_p0),
    .din1(wgt_M_instance_6_V_reg_5396),
    .dout(mul_ln1352_6_fu_2802_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U9(
    .din0(mul_ln1352_7_fu_2829_p0),
    .din1(wgt_M_instance_7_V_reg_5401),
    .dout(mul_ln1352_7_fu_2829_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U10(
    .din0(mul_ln1352_8_fu_2866_p0),
    .din1(wgt_M_instance_0_V_1_reg_5406),
    .dout(mul_ln1352_8_fu_2866_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U11(
    .din0(mul_ln1352_9_fu_2879_p0),
    .din1(wgt_M_instance_1_V_1_reg_5411),
    .dout(mul_ln1352_9_fu_2879_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U12(
    .din0(mul_ln1352_10_fu_2892_p0),
    .din1(wgt_M_instance_2_V_1_reg_5416),
    .dout(mul_ln1352_10_fu_2892_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U13(
    .din0(mul_ln1352_11_fu_2905_p0),
    .din1(wgt_M_instance_3_V_1_reg_5421),
    .dout(mul_ln1352_11_fu_2905_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U14(
    .din0(mul_ln1352_12_fu_2918_p0),
    .din1(wgt_M_instance_4_V_1_reg_5426),
    .dout(mul_ln1352_12_fu_2918_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U15(
    .din0(mul_ln1352_13_fu_2931_p0),
    .din1(wgt_M_instance_5_V_1_reg_5431),
    .dout(mul_ln1352_13_fu_2931_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U16(
    .din0(mul_ln1352_14_fu_2940_p0),
    .din1(wgt_M_instance_6_V_1_reg_5436),
    .dout(mul_ln1352_14_fu_2940_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U17(
    .din0(mul_ln1352_15_fu_2953_p0),
    .din1(wgt_M_instance_7_V_1_reg_5441),
    .dout(mul_ln1352_15_fu_2953_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U18(
    .din0(mul_ln1352_16_fu_2990_p0),
    .din1(wgt_M_instance_0_V_2_reg_5446),
    .dout(mul_ln1352_16_fu_2990_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U19(
    .din0(mul_ln1352_17_fu_3003_p0),
    .din1(wgt_M_instance_1_V_2_reg_5451),
    .dout(mul_ln1352_17_fu_3003_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U20(
    .din0(mul_ln1352_18_fu_3016_p0),
    .din1(wgt_M_instance_2_V_2_reg_5456),
    .dout(mul_ln1352_18_fu_3016_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U21(
    .din0(mul_ln1352_19_fu_3029_p0),
    .din1(wgt_M_instance_3_V_2_reg_5461),
    .dout(mul_ln1352_19_fu_3029_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U22(
    .din0(mul_ln1352_20_fu_3042_p0),
    .din1(wgt_M_instance_4_V_2_reg_5466),
    .dout(mul_ln1352_20_fu_3042_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U23(
    .din0(mul_ln1352_21_fu_3055_p0),
    .din1(wgt_M_instance_5_V_2_reg_5471),
    .dout(mul_ln1352_21_fu_3055_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U24(
    .din0(mul_ln1352_22_fu_3064_p0),
    .din1(wgt_M_instance_6_V_2_reg_5476),
    .dout(mul_ln1352_22_fu_3064_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U25(
    .din0(mul_ln1352_23_fu_3077_p0),
    .din1(wgt_M_instance_7_V_2_reg_5481),
    .dout(mul_ln1352_23_fu_3077_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U26(
    .din0(mul_ln1352_24_fu_3114_p0),
    .din1(wgt_M_instance_0_V_3_reg_5486),
    .dout(mul_ln1352_24_fu_3114_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U27(
    .din0(mul_ln1352_25_fu_3127_p0),
    .din1(wgt_M_instance_1_V_3_reg_5491),
    .dout(mul_ln1352_25_fu_3127_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U28(
    .din0(mul_ln1352_26_fu_3140_p0),
    .din1(wgt_M_instance_2_V_3_reg_5496),
    .dout(mul_ln1352_26_fu_3140_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U29(
    .din0(mul_ln1352_27_fu_3153_p0),
    .din1(wgt_M_instance_3_V_3_reg_5501),
    .dout(mul_ln1352_27_fu_3153_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U30(
    .din0(mul_ln1352_28_fu_3166_p0),
    .din1(wgt_M_instance_4_V_3_reg_5506),
    .dout(mul_ln1352_28_fu_3166_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U31(
    .din0(mul_ln1352_29_fu_3179_p0),
    .din1(wgt_M_instance_5_V_3_reg_5511),
    .dout(mul_ln1352_29_fu_3179_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U32(
    .din0(mul_ln1352_30_fu_3188_p0),
    .din1(wgt_M_instance_6_V_3_reg_5516),
    .dout(mul_ln1352_30_fu_3188_p2)
);

StreamingFCLayer_Batch_4_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U33(
    .din0(mul_ln1352_31_fu_3201_p0),
    .din1(wgt_M_instance_7_V_3_reg_5521),
    .dout(mul_ln1352_31_fu_3201_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd0) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470 <= inElem_V_1_fu_1835_p66;
    end else if ((((trunc_ln321_fu_1969_p1 == 6'd46) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd47) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd48) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd49) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd50) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd51) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd52) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd53) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd54) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd55) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd56) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd57) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd58) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd59) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd60) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd61) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd62) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd63) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd2) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd3) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd4) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd5) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd6) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd7) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd8) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd9) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd10) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd11) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd12) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd13) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd14) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd15) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd16) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd17) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd18) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd19) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd20) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd21) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd22) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd23) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd24) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd25) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd26) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd27) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd28) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd29) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd30) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd31) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd32) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd33) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd34) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd35) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd36) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd37) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd38) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd39) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd40) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd41) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd42) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd43) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd44) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_1969_p1 == 6'd45) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470 <= in_V_V_TDATA;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470 <= ap_phi_reg_pp0_iter0_act_m_val_V_reg_1470;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_reg_1459 <= i_fu_1621_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_reg_1459 <= 14'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_5526 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        nf_assign_fu_708 <= select_ln301_fu_3310_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        nf_assign_fu_708 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_2622_p2 == 1'd0) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        sf_1_fu_448 <= sf_fu_2616_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_2622_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        sf_1_fu_448 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        accu_V_0_0_0_fu_432 <= accu_0_0_V_fu_3397_p2;
        accu_V_0_1_0_fu_436 <= accu_0_1_V_fu_3437_p2;
        accu_V_0_2_0_fu_440 <= accu_0_2_V_fu_3477_p2;
        accu_V_0_3_0_fu_444 <= accu_0_3_V_fu_3517_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln700_11_reg_5560 <= add_ln700_11_fu_2969_p2;
        add_ln700_13_reg_5565 <= add_ln700_13_fu_2981_p2;
        add_ln700_17_reg_5575 <= add_ln700_17_fu_3087_p2;
        add_ln700_19_reg_5580 <= add_ln700_19_fu_3093_p2;
        add_ln700_1_reg_5535 <= add_ln700_1_fu_2839_p2;
        add_ln700_21_reg_5585 <= add_ln700_21_fu_3105_p2;
        add_ln700_25_reg_5595 <= add_ln700_25_fu_3211_p2;
        add_ln700_27_reg_5600 <= add_ln700_27_fu_3217_p2;
        add_ln700_29_reg_5605 <= add_ln700_29_fu_3229_p2;
        add_ln700_3_reg_5540 <= add_ln700_3_fu_2845_p2;
        add_ln700_5_reg_5545 <= add_ln700_5_fu_2857_p2;
        add_ln700_9_reg_5555 <= add_ln700_9_fu_2963_p2;
        icmp_ln271_reg_5358_pp0_iter1_reg <= icmp_ln271_reg_5358;
        icmp_ln289_reg_5526_pp0_iter1_reg <= icmp_ln289_reg_5526;
        mul_ln1352_13_reg_5550 <= mul_ln1352_13_fu_2931_p2;
        mul_ln1352_21_reg_5570 <= mul_ln1352_21_fu_3055_p2;
        mul_ln1352_29_reg_5590 <= mul_ln1352_29_fu_3179_p2;
        mul_ln1352_5_reg_5530 <= mul_ln1352_5_fu_2779_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_5526_pp0_iter2_reg == 1'd1))) begin
        add_ln700_36_reg_6170 <= add_ln700_36_fu_3998_p2;
        add_ln700_43_reg_6175 <= add_ln700_43_fu_4046_p2;
        add_ln700_49_reg_6180 <= add_ln700_49_fu_4171_p2;
        add_ln700_56_reg_6185 <= add_ln700_56_fu_4219_p2;
        add_ln700_62_reg_6190 <= add_ln700_62_fu_4344_p2;
        add_ln700_69_reg_6195 <= add_ln700_69_fu_4392_p2;
        add_ln700_75_reg_6200 <= add_ln700_75_fu_4517_p2;
        add_ln700_82_reg_6205 <= add_ln700_82_fu_4565_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_1615_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln271_reg_5358 <= icmp_ln271_fu_2296_p2;
        icmp_ln289_reg_5526 <= icmp_ln289_fu_2622_p2;
        wgt_M_instance_0_V_1_reg_5406 <= {{weight_V_V_TDATA[35:32]}};
        wgt_M_instance_0_V_2_reg_5446 <= {{weight_V_V_TDATA[67:64]}};
        wgt_M_instance_0_V_3_reg_5486 <= {{weight_V_V_TDATA[99:96]}};
        wgt_M_instance_0_V_reg_5366 <= wgt_M_instance_0_V_fu_2302_p1;
        wgt_M_instance_1_V_1_reg_5411 <= {{weight_V_V_TDATA[39:36]}};
        wgt_M_instance_1_V_2_reg_5451 <= {{weight_V_V_TDATA[71:68]}};
        wgt_M_instance_1_V_3_reg_5491 <= {{weight_V_V_TDATA[103:100]}};
        wgt_M_instance_1_V_reg_5371 <= {{weight_V_V_TDATA[7:4]}};
        wgt_M_instance_2_V_1_reg_5416 <= {{weight_V_V_TDATA[43:40]}};
        wgt_M_instance_2_V_2_reg_5456 <= {{weight_V_V_TDATA[75:72]}};
        wgt_M_instance_2_V_3_reg_5496 <= {{weight_V_V_TDATA[107:104]}};
        wgt_M_instance_2_V_reg_5376 <= {{weight_V_V_TDATA[11:8]}};
        wgt_M_instance_3_V_1_reg_5421 <= {{weight_V_V_TDATA[47:44]}};
        wgt_M_instance_3_V_2_reg_5461 <= {{weight_V_V_TDATA[79:76]}};
        wgt_M_instance_3_V_3_reg_5501 <= {{weight_V_V_TDATA[111:108]}};
        wgt_M_instance_3_V_reg_5381 <= {{weight_V_V_TDATA[15:12]}};
        wgt_M_instance_4_V_1_reg_5426 <= {{weight_V_V_TDATA[51:48]}};
        wgt_M_instance_4_V_2_reg_5466 <= {{weight_V_V_TDATA[83:80]}};
        wgt_M_instance_4_V_3_reg_5506 <= {{weight_V_V_TDATA[115:112]}};
        wgt_M_instance_4_V_reg_5386 <= {{weight_V_V_TDATA[19:16]}};
        wgt_M_instance_5_V_1_reg_5431 <= {{weight_V_V_TDATA[55:52]}};
        wgt_M_instance_5_V_2_reg_5471 <= {{weight_V_V_TDATA[87:84]}};
        wgt_M_instance_5_V_3_reg_5511 <= {{weight_V_V_TDATA[119:116]}};
        wgt_M_instance_5_V_reg_5391 <= {{weight_V_V_TDATA[23:20]}};
        wgt_M_instance_6_V_1_reg_5436 <= {{weight_V_V_TDATA[59:56]}};
        wgt_M_instance_6_V_2_reg_5476 <= {{weight_V_V_TDATA[91:88]}};
        wgt_M_instance_6_V_3_reg_5516 <= {{weight_V_V_TDATA[123:120]}};
        wgt_M_instance_6_V_reg_5396 <= {{weight_V_V_TDATA[27:24]}};
        wgt_M_instance_7_V_1_reg_5441 <= {{weight_V_V_TDATA[63:60]}};
        wgt_M_instance_7_V_2_reg_5481 <= {{weight_V_V_TDATA[95:92]}};
        wgt_M_instance_7_V_3_reg_5521 <= {{weight_V_V_TDATA[127:124]}};
        wgt_M_instance_7_V_reg_5401 <= {{weight_V_V_TDATA[31:28]}};
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln289_reg_5526_pp0_iter2_reg <= icmp_ln289_reg_5526_pp0_iter1_reg;
        icmp_ln289_reg_5526_pp0_iter3_reg <= icmp_ln289_reg_5526_pp0_iter2_reg;
        icmp_ln899_14_reg_5960_pp0_iter3_reg <= icmp_ln899_14_reg_5960;
        icmp_ln899_15_reg_5965_pp0_iter3_reg <= icmp_ln899_15_reg_5965;
        icmp_ln899_16_reg_5970_pp0_iter3_reg <= icmp_ln899_16_reg_5970;
        icmp_ln899_1_reg_5895_pp0_iter3_reg <= icmp_ln899_1_reg_5895;
        icmp_ln899_28_reg_6030_pp0_iter3_reg <= icmp_ln899_28_reg_6030;
        icmp_ln899_29_reg_6035_pp0_iter3_reg <= icmp_ln899_29_reg_6035;
        icmp_ln899_2_reg_5900_pp0_iter3_reg <= icmp_ln899_2_reg_5900;
        icmp_ln899_30_reg_6040_pp0_iter3_reg <= icmp_ln899_30_reg_6040;
        icmp_ln899_42_reg_6100_pp0_iter3_reg <= icmp_ln899_42_reg_6100;
        icmp_ln899_43_reg_6105_pp0_iter3_reg <= icmp_ln899_43_reg_6105;
        icmp_ln899_44_reg_6110_pp0_iter3_reg <= icmp_ln899_44_reg_6110;
        icmp_ln899_reg_5890_pp0_iter3_reg <= icmp_ln899_reg_5890;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_5526_pp0_iter1_reg == 1'd1))) begin
        icmp_ln899_10_reg_5940 <= icmp_ln899_10_fu_3603_p2;
        icmp_ln899_11_reg_5945 <= icmp_ln899_11_fu_3609_p2;
        icmp_ln899_12_reg_5950 <= icmp_ln899_12_fu_3615_p2;
        icmp_ln899_13_reg_5955 <= icmp_ln899_13_fu_3621_p2;
        icmp_ln899_14_reg_5960 <= icmp_ln899_14_fu_3627_p2;
        icmp_ln899_15_reg_5965 <= icmp_ln899_15_fu_3633_p2;
        icmp_ln899_16_reg_5970 <= icmp_ln899_16_fu_3639_p2;
        icmp_ln899_17_reg_5975 <= icmp_ln899_17_fu_3645_p2;
        icmp_ln899_18_reg_5980 <= icmp_ln899_18_fu_3651_p2;
        icmp_ln899_19_reg_5985 <= icmp_ln899_19_fu_3657_p2;
        icmp_ln899_1_reg_5895 <= icmp_ln899_1_fu_3549_p2;
        icmp_ln899_20_reg_5990 <= icmp_ln899_20_fu_3663_p2;
        icmp_ln899_21_reg_5995 <= icmp_ln899_21_fu_3669_p2;
        icmp_ln899_22_reg_6000 <= icmp_ln899_22_fu_3675_p2;
        icmp_ln899_23_reg_6005 <= icmp_ln899_23_fu_3681_p2;
        icmp_ln899_24_reg_6010 <= icmp_ln899_24_fu_3687_p2;
        icmp_ln899_25_reg_6015 <= icmp_ln899_25_fu_3693_p2;
        icmp_ln899_26_reg_6020 <= icmp_ln899_26_fu_3699_p2;
        icmp_ln899_27_reg_6025 <= icmp_ln899_27_fu_3705_p2;
        icmp_ln899_28_reg_6030 <= icmp_ln899_28_fu_3711_p2;
        icmp_ln899_29_reg_6035 <= icmp_ln899_29_fu_3717_p2;
        icmp_ln899_2_reg_5900 <= icmp_ln899_2_fu_3555_p2;
        icmp_ln899_30_reg_6040 <= icmp_ln899_30_fu_3723_p2;
        icmp_ln899_31_reg_6045 <= icmp_ln899_31_fu_3729_p2;
        icmp_ln899_32_reg_6050 <= icmp_ln899_32_fu_3735_p2;
        icmp_ln899_33_reg_6055 <= icmp_ln899_33_fu_3741_p2;
        icmp_ln899_34_reg_6060 <= icmp_ln899_34_fu_3747_p2;
        icmp_ln899_35_reg_6065 <= icmp_ln899_35_fu_3753_p2;
        icmp_ln899_36_reg_6070 <= icmp_ln899_36_fu_3759_p2;
        icmp_ln899_37_reg_6075 <= icmp_ln899_37_fu_3765_p2;
        icmp_ln899_38_reg_6080 <= icmp_ln899_38_fu_3771_p2;
        icmp_ln899_39_reg_6085 <= icmp_ln899_39_fu_3777_p2;
        icmp_ln899_3_reg_5905 <= icmp_ln899_3_fu_3561_p2;
        icmp_ln899_40_reg_6090 <= icmp_ln899_40_fu_3783_p2;
        icmp_ln899_41_reg_6095 <= icmp_ln899_41_fu_3789_p2;
        icmp_ln899_42_reg_6100 <= icmp_ln899_42_fu_3795_p2;
        icmp_ln899_43_reg_6105 <= icmp_ln899_43_fu_3801_p2;
        icmp_ln899_44_reg_6110 <= icmp_ln899_44_fu_3807_p2;
        icmp_ln899_45_reg_6115 <= icmp_ln899_45_fu_3813_p2;
        icmp_ln899_46_reg_6120 <= icmp_ln899_46_fu_3819_p2;
        icmp_ln899_47_reg_6125 <= icmp_ln899_47_fu_3825_p2;
        icmp_ln899_48_reg_6130 <= icmp_ln899_48_fu_3831_p2;
        icmp_ln899_49_reg_6135 <= icmp_ln899_49_fu_3837_p2;
        icmp_ln899_4_reg_5910 <= icmp_ln899_4_fu_3567_p2;
        icmp_ln899_50_reg_6140 <= icmp_ln899_50_fu_3843_p2;
        icmp_ln899_51_reg_6145 <= icmp_ln899_51_fu_3849_p2;
        icmp_ln899_52_reg_6150 <= icmp_ln899_52_fu_3855_p2;
        icmp_ln899_53_reg_6155 <= icmp_ln899_53_fu_3861_p2;
        icmp_ln899_54_reg_6160 <= icmp_ln899_54_fu_3867_p2;
        icmp_ln899_55_reg_6165 <= icmp_ln899_55_fu_3873_p2;
        icmp_ln899_5_reg_5915 <= icmp_ln899_5_fu_3573_p2;
        icmp_ln899_6_reg_5920 <= icmp_ln899_6_fu_3579_p2;
        icmp_ln899_7_reg_5925 <= icmp_ln899_7_fu_3585_p2;
        icmp_ln899_8_reg_5930 <= icmp_ln899_8_fu_3591_p2;
        icmp_ln899_9_reg_5935 <= icmp_ln899_9_fu_3597_p2;
        icmp_ln899_reg_5890 <= icmp_ln899_fu_3543_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd9) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_10_fu_488 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd10) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_11_fu_492 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd11) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_12_fu_496 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd12) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_13_fu_500 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd13) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_14_fu_504 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd14) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_15_fu_508 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd15) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_16_fu_512 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd16) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_17_fu_516 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd17) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_18_fu_520 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd18) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_19_fu_524 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_1_fu_456 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd19) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_20_fu_528 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd20) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_21_fu_532 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd21) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_22_fu_536 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd22) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_23_fu_540 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd23) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_24_fu_544 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd24) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_25_fu_548 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd25) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_26_fu_552 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd26) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_27_fu_556 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd27) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_28_fu_560 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd28) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_29_fu_564 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd2) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_2_fu_460 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd29) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_30_fu_568 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd30) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_31_fu_572 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd31) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_32_fu_576 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd32) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_33_fu_580 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd33) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_34_fu_584 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd34) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_35_fu_588 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd35) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_36_fu_592 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd36) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_37_fu_596 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd37) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_38_fu_600 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd38) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_39_fu_604 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd39) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_40_fu_608 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd40) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_41_fu_612 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd41) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_42_fu_616 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd42) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_43_fu_620 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd43) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_44_fu_624 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd44) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_45_fu_628 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd45) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_46_fu_632 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd46) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_47_fu_636 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd47) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_48_fu_640 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd48) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_49_fu_644 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd3) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_4_fu_464 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd49) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_50_fu_648 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd50) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_51_fu_652 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd51) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_52_fu_656 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd52) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_53_fu_660 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd53) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_54_fu_664 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd54) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_55_fu_668 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd55) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_56_fu_672 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd56) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_57_fu_676 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd57) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_58_fu_680 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd58) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_59_fu_684 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd4) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_5_fu_468 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd59) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_60_fu_688 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd60) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_61_fu_692 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd61) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_62_fu_696 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd62) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_63_fu_700 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd63) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_64_fu_704 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd5) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_6_fu_472 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd6) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_7_fu_476 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd7) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_8_fu_480 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd8) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_9_fu_484 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_1969_p1 == 6'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_fu_452 <= in_V_V_TDATA;
    end
end

always @ (*) begin
    if ((icmp_ln248_fu_1615_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state7) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_5526 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_sig_allocacmp_nf_assign_load_1 = select_ln301_fu_3310_p3;
    end else begin
        ap_sig_allocacmp_nf_assign_load_1 = nf_assign_fu_708;
    end
end

always @ (*) begin
    if (((icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op162_read_state2 == 1'b1))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_5526_pp0_iter3_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_5526_pp0_iter3_reg == 1'd1) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_10_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_10_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_11_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_11_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_12_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_12_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_13_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_13_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_14_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_14_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_15_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_15_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_16_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_16_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_17_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_17_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_18_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_18_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_19_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_19_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_1_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_1_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_20_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_20_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_21_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_21_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_22_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_22_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_23_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_23_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_24_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_24_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_25_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_25_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_26_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_26_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_27_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_27_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_28_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_28_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_29_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_29_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_2_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_2_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_30_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_30_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_31_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_31_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_32_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_32_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_33_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_33_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_34_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_34_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_35_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_35_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_36_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_36_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_37_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_37_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_38_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_38_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_39_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_39_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_3_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_3_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_40_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_40_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_41_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_41_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_42_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_42_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_43_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_43_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_44_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_44_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_45_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_45_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_46_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_46_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_47_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_47_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_48_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_48_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_49_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_49_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_4_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_4_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_50_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_50_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_51_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_51_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_52_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_52_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_53_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_53_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_54_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_54_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_55_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_55_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_5_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_5_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_6_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_6_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_7_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_7_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_8_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_8_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_9_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_9_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln248_fu_1615_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TDATA_blk_n = weight_V_V_TVALID;
    end else begin
        weight_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_1615_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TREADY = 1'b1;
    end else begin
        weight_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln248_fu_1615_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((ap_enable_reg_pp0_iter3 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter3 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln248_fu_1615_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accu_0_0_V_fu_3397_p2 = ($signed(add_ln700_2_fu_3375_p2) + $signed(sext_ln700_5_fu_3393_p1));

assign accu_0_1_V_fu_3437_p2 = ($signed(add_ln700_10_fu_3415_p2) + $signed(sext_ln700_11_fu_3433_p1));

assign accu_0_2_V_fu_3477_p2 = ($signed(add_ln700_18_fu_3455_p2) + $signed(sext_ln700_17_fu_3473_p1));

assign accu_0_3_V_fu_3517_p2 = ($signed(add_ln700_26_fu_3495_p2) + $signed(sext_ln700_23_fu_3513_p1));

assign add_ln700_10_fu_3415_p2 = ($signed(add_ln700_8_fu_3406_p2) + $signed(sext_ln700_8_fu_3412_p1));

assign add_ln700_11_fu_2969_p2 = ($signed(sext_ln170_6_fu_2872_p1) + $signed(sext_ln170_9_fu_2911_p1));

assign add_ln700_12_fu_2975_p2 = ($signed(sext_ln700_7_fu_2959_p1) + $signed(sext_ln170_7_fu_2885_p1));

assign add_ln700_13_fu_2981_p2 = ($signed(sext_ln170_8_fu_2898_p1) + $signed(add_ln700_12_fu_2975_p2));

assign add_ln700_14_fu_3427_p2 = ($signed(sext_ln700_9_fu_3421_p1) + $signed(sext_ln700_10_fu_3424_p1));

assign add_ln700_16_fu_3446_p2 = ($signed(sext_ln700_12_fu_3443_p1) + $signed(select_ln271_1_fu_3342_p3));

assign add_ln700_17_fu_3087_p2 = ($signed(sext_ln170_16_fu_3048_p1) + $signed(sext_ln170_17_fu_3070_p1));

assign add_ln700_18_fu_3455_p2 = ($signed(add_ln700_16_fu_3446_p2) + $signed(sext_ln700_14_fu_3452_p1));

assign add_ln700_19_fu_3093_p2 = ($signed(sext_ln170_12_fu_2996_p1) + $signed(sext_ln170_15_fu_3035_p1));

assign add_ln700_1_fu_2839_p2 = ($signed(sext_ln170_4_fu_2758_p1) + $signed(sext_ln170_5_fu_2808_p1));

assign add_ln700_20_fu_3099_p2 = ($signed(sext_ln700_13_fu_3083_p1) + $signed(sext_ln170_13_fu_3009_p1));

assign add_ln700_21_fu_3105_p2 = ($signed(sext_ln170_14_fu_3022_p1) + $signed(add_ln700_20_fu_3099_p2));

assign add_ln700_22_fu_3467_p2 = ($signed(sext_ln700_15_fu_3461_p1) + $signed(sext_ln700_16_fu_3464_p1));

assign add_ln700_24_fu_3486_p2 = ($signed(sext_ln700_18_fu_3483_p1) + $signed(select_ln271_fu_3335_p3));

assign add_ln700_25_fu_3211_p2 = ($signed(sext_ln170_22_fu_3172_p1) + $signed(sext_ln170_23_fu_3194_p1));

assign add_ln700_26_fu_3495_p2 = ($signed(add_ln700_24_fu_3486_p2) + $signed(sext_ln700_20_fu_3492_p1));

assign add_ln700_27_fu_3217_p2 = ($signed(sext_ln170_18_fu_3120_p1) + $signed(sext_ln170_21_fu_3159_p1));

assign add_ln700_28_fu_3223_p2 = ($signed(sext_ln700_19_fu_3207_p1) + $signed(sext_ln170_19_fu_3133_p1));

assign add_ln700_29_fu_3229_p2 = ($signed(sext_ln170_20_fu_3146_p1) + $signed(add_ln700_28_fu_3223_p2));

assign add_ln700_2_fu_3375_p2 = ($signed(add_ln700_fu_3366_p2) + $signed(sext_ln700_2_fu_3372_p1));

assign add_ln700_30_fu_3507_p2 = ($signed(sext_ln700_21_fu_3501_p1) + $signed(sext_ln700_22_fu_3504_p1));

assign add_ln700_32_fu_4602_p2 = (zext_ln142_1_fu_4589_p1 + zext_ln142_2_fu_4598_p1);

assign add_ln700_33_fu_4612_p2 = (zext_ln700_1_fu_4608_p1 + select_ln700_fu_4576_p3);

assign add_ln700_34_fu_3978_p2 = (zext_ln142_3_fu_3884_p1 + zext_ln142_4_fu_3893_p1);

assign add_ln700_35_fu_3988_p2 = (zext_ln142_5_fu_3902_p1 + zext_ln142_6_fu_3911_p1);

assign add_ln700_36_fu_3998_p2 = (zext_ln700_3_fu_3994_p1 + zext_ln700_2_fu_3984_p1);

assign add_ln700_37_fu_4621_p2 = (zext_ln700_4_fu_4618_p1 + add_ln700_33_fu_4612_p2);

assign add_ln700_38_fu_4004_p2 = (zext_ln142_8_fu_3929_p1 + zext_ln142_9_fu_3938_p1);

assign add_ln700_39_fu_4010_p2 = (add_ln700_38_fu_4004_p2 + zext_ln142_7_fu_3920_p1);

assign add_ln700_3_fu_2845_p2 = ($signed(sext_ln170_fu_2650_p1) + $signed(sext_ln170_3_fu_2731_p1));

assign add_ln700_40_fu_4020_p2 = (zext_ln142_10_fu_3947_p1 + zext_ln142_11_fu_3956_p1);

assign add_ln700_41_fu_4030_p2 = (zext_ln142_12_fu_3965_p1 + zext_ln700_fu_3974_p1);

assign add_ln700_42_fu_4040_p2 = (zext_ln700_7_fu_4036_p1 + zext_ln700_6_fu_4026_p1);

assign add_ln700_43_fu_4046_p2 = (add_ln700_42_fu_4040_p2 + zext_ln700_5_fu_4016_p1);

assign add_ln700_44_fu_4630_p2 = (zext_ln700_8_fu_4627_p1 + add_ln700_37_fu_4621_p2);

assign add_ln700_45_fu_4667_p2 = (zext_ln142_13_fu_4654_p1 + zext_ln142_14_fu_4663_p1);

assign add_ln700_46_fu_4677_p2 = (zext_ln700_10_fu_4673_p1 + select_ln700_1_fu_4641_p3);

assign add_ln700_47_fu_4151_p2 = (zext_ln142_15_fu_4057_p1 + zext_ln142_16_fu_4066_p1);

assign add_ln700_48_fu_4161_p2 = (zext_ln142_17_fu_4075_p1 + zext_ln142_18_fu_4084_p1);

assign add_ln700_49_fu_4171_p2 = (zext_ln700_12_fu_4167_p1 + zext_ln700_11_fu_4157_p1);

assign add_ln700_4_fu_2851_p2 = ($signed(sext_ln700_1_fu_2835_p1) + $signed(sext_ln170_1_fu_2677_p1));

assign add_ln700_50_fu_4686_p2 = (zext_ln700_13_fu_4683_p1 + add_ln700_46_fu_4677_p2);

assign add_ln700_51_fu_4177_p2 = (zext_ln142_20_fu_4102_p1 + zext_ln142_21_fu_4111_p1);

assign add_ln700_52_fu_4183_p2 = (add_ln700_51_fu_4177_p2 + zext_ln142_19_fu_4093_p1);

assign add_ln700_53_fu_4193_p2 = (zext_ln142_22_fu_4120_p1 + zext_ln142_23_fu_4129_p1);

assign add_ln700_54_fu_4203_p2 = (zext_ln142_24_fu_4138_p1 + zext_ln700_9_fu_4147_p1);

assign add_ln700_55_fu_4213_p2 = (zext_ln700_16_fu_4209_p1 + zext_ln700_15_fu_4199_p1);

assign add_ln700_56_fu_4219_p2 = (add_ln700_55_fu_4213_p2 + zext_ln700_14_fu_4189_p1);

assign add_ln700_57_fu_4695_p2 = (zext_ln700_17_fu_4692_p1 + add_ln700_50_fu_4686_p2);

assign add_ln700_58_fu_4732_p2 = (zext_ln142_25_fu_4719_p1 + zext_ln142_26_fu_4728_p1);

assign add_ln700_59_fu_4742_p2 = (zext_ln700_19_fu_4738_p1 + select_ln700_2_fu_4706_p3);

assign add_ln700_5_fu_2857_p2 = ($signed(sext_ln170_2_fu_2704_p1) + $signed(add_ln700_4_fu_2851_p2));

assign add_ln700_60_fu_4324_p2 = (zext_ln142_27_fu_4230_p1 + zext_ln142_28_fu_4239_p1);

assign add_ln700_61_fu_4334_p2 = (zext_ln142_29_fu_4248_p1 + zext_ln142_30_fu_4257_p1);

assign add_ln700_62_fu_4344_p2 = (zext_ln700_21_fu_4340_p1 + zext_ln700_20_fu_4330_p1);

assign add_ln700_63_fu_4751_p2 = (zext_ln700_22_fu_4748_p1 + add_ln700_59_fu_4742_p2);

assign add_ln700_64_fu_4350_p2 = (zext_ln142_32_fu_4275_p1 + zext_ln142_33_fu_4284_p1);

assign add_ln700_65_fu_4356_p2 = (add_ln700_64_fu_4350_p2 + zext_ln142_31_fu_4266_p1);

assign add_ln700_66_fu_4366_p2 = (zext_ln142_34_fu_4293_p1 + zext_ln142_35_fu_4302_p1);

assign add_ln700_67_fu_4376_p2 = (zext_ln142_36_fu_4311_p1 + zext_ln700_18_fu_4320_p1);

assign add_ln700_68_fu_4386_p2 = (zext_ln700_25_fu_4382_p1 + zext_ln700_24_fu_4372_p1);

assign add_ln700_69_fu_4392_p2 = (add_ln700_68_fu_4386_p2 + zext_ln700_23_fu_4362_p1);

assign add_ln700_6_fu_3387_p2 = ($signed(sext_ln700_3_fu_3381_p1) + $signed(sext_ln700_4_fu_3384_p1));

assign add_ln700_70_fu_4760_p2 = (zext_ln700_26_fu_4757_p1 + add_ln700_63_fu_4751_p2);

assign add_ln700_71_fu_4797_p2 = (zext_ln142_37_fu_4784_p1 + zext_ln142_38_fu_4793_p1);

assign add_ln700_72_fu_4807_p2 = (zext_ln700_28_fu_4803_p1 + select_ln700_3_fu_4771_p3);

assign add_ln700_73_fu_4497_p2 = (zext_ln142_39_fu_4403_p1 + zext_ln142_40_fu_4412_p1);

assign add_ln700_74_fu_4507_p2 = (zext_ln142_41_fu_4421_p1 + zext_ln142_42_fu_4430_p1);

assign add_ln700_75_fu_4517_p2 = (zext_ln700_30_fu_4513_p1 + zext_ln700_29_fu_4503_p1);

assign add_ln700_76_fu_4816_p2 = (zext_ln700_31_fu_4813_p1 + add_ln700_72_fu_4807_p2);

assign add_ln700_77_fu_4523_p2 = (zext_ln142_44_fu_4448_p1 + zext_ln142_45_fu_4457_p1);

assign add_ln700_78_fu_4529_p2 = (add_ln700_77_fu_4523_p2 + zext_ln142_43_fu_4439_p1);

assign add_ln700_79_fu_4539_p2 = (zext_ln142_46_fu_4466_p1 + zext_ln142_47_fu_4475_p1);

assign add_ln700_80_fu_4549_p2 = (zext_ln142_48_fu_4484_p1 + zext_ln700_27_fu_4493_p1);

assign add_ln700_81_fu_4559_p2 = (zext_ln700_34_fu_4555_p1 + zext_ln700_33_fu_4545_p1);

assign add_ln700_82_fu_4565_p2 = (add_ln700_81_fu_4559_p2 + zext_ln700_32_fu_4535_p1);

assign add_ln700_83_fu_4825_p2 = (zext_ln700_35_fu_4822_p1 + add_ln700_76_fu_4816_p2);

assign add_ln700_8_fu_3406_p2 = ($signed(sext_ln700_6_fu_3403_p1) + $signed(select_ln271_2_fu_3349_p3));

assign add_ln700_9_fu_2963_p2 = ($signed(sext_ln170_10_fu_2924_p1) + $signed(sext_ln170_11_fu_2946_p1));

assign add_ln700_fu_3366_p2 = ($signed(sext_ln700_fu_3363_p1) + $signed(select_ln271_3_fu_3356_p3));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((icmp_ln248_fu_1615_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_block_state6_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((icmp_ln248_fu_1615_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_block_state6_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((icmp_ln248_fu_1615_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op162_read_state2 == 1'b1)) | ((icmp_ln248_fu_1615_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state6_io = ((icmp_ln289_reg_5526_pp0_iter3_reg == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_reg_pp0_iter0_act_m_val_V_reg_1470 = 'bx;

always @ (*) begin
    ap_predicate_op162_read_state2 = ((icmp_ln252_fu_1630_p2 == 1'd1) & (icmp_ln248_fu_1615_p2 == 1'd0));
end

assign arg_V_read_assign_1_fu_2654_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470[7:4]}};

assign arg_V_read_assign_2_fu_2681_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470[11:8]}};

assign arg_V_read_assign_3_fu_2708_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470[15:12]}};

assign arg_V_read_assign_4_fu_2735_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470[19:16]}};

assign arg_V_read_assign_5_fu_2762_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470[23:20]}};

assign arg_V_read_assign_6_fu_2785_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470[27:24]}};

assign arg_V_read_assign_7_fu_2812_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470[31:28]}};

assign i_fu_1621_p2 = (i_0_reg_1459 + 14'd1);

assign icmp_ln248_fu_1615_p2 = ((i_0_reg_1459 == 14'd8192) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_1630_p2 = ((ap_sig_allocacmp_nf_assign_load_1 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln271_fu_2296_p2 = ((sf_1_fu_448 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln289_fu_2622_p2 = ((sf_fu_2616_p2 == 32'd64) ? 1'b1 : 1'b0);

assign icmp_ln301_fu_3304_p2 = ((nf_fu_3298_p2 == 32'd128) ? 1'b1 : 1'b0);

assign icmp_ln899_10_fu_3603_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_53_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_11_fu_3609_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_52_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_12_fu_3615_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_51_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_13_fu_3621_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_50_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_14_fu_3627_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_41_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_15_fu_3633_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_40_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_16_fu_3639_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_35_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_17_fu_3645_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_34_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_18_fu_3651_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_33_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_19_fu_3657_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_32_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_1_fu_3549_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_54_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_20_fu_3663_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_31_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_21_fu_3669_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_30_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_22_fu_3675_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_29_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_23_fu_3681_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_28_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_24_fu_3687_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_39_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_25_fu_3693_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_38_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_26_fu_3699_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_37_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_27_fu_3705_p2 = (($signed(accu_0_1_V_fu_3437_p2) < $signed(threshs_m_thresholds_36_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_28_fu_3711_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_27_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_29_fu_3717_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_26_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_2_fu_3555_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_49_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_30_fu_3723_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_21_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_31_fu_3729_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_20_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_32_fu_3735_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_19_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_33_fu_3741_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_18_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_34_fu_3747_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_17_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_35_fu_3753_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_16_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_36_fu_3759_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_15_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_37_fu_3765_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_14_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_38_fu_3771_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_25_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_39_fu_3777_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_24_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_3_fu_3561_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_48_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_40_fu_3783_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_23_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_41_fu_3789_p2 = (($signed(accu_0_2_V_fu_3477_p2) < $signed(threshs_m_thresholds_22_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_42_fu_3795_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_13_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_43_fu_3801_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_12_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_44_fu_3807_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_7_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_45_fu_3813_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_6_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_46_fu_3819_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_5_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_47_fu_3825_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_4_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_48_fu_3831_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_3_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_49_fu_3837_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_2_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_4_fu_3567_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_47_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_50_fu_3843_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_1_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_51_fu_3849_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_52_fu_3855_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_11_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_53_fu_3861_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_10_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_54_fu_3867_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_9_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_55_fu_3873_p2 = (($signed(accu_0_3_V_fu_3517_p2) < $signed(threshs_m_thresholds_8_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_5_fu_3573_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_46_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_6_fu_3579_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_45_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_7_fu_3585_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_44_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_8_fu_3591_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_43_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_9_fu_3597_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_42_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_fu_3543_p2 = (($signed(accu_0_0_V_fu_3397_p2) < $signed(threshs_m_thresholds_55_q0)) ? 1'b1 : 1'b0);

assign inElem_V_1_fu_1835_p65 = sf_1_fu_448[5:0];

assign mul_ln1352_10_fu_2892_p0 = sext_ln215_5_fu_2694_p1;

assign mul_ln1352_11_fu_2905_p0 = sext_ln215_7_fu_2721_p1;

assign mul_ln1352_12_fu_2918_p0 = sext_ln215_9_fu_2748_p1;

assign mul_ln1352_13_fu_2931_p0 = sext_ln215_11_fu_2775_p1;

assign mul_ln1352_14_fu_2940_p0 = sext_ln215_13_fu_2798_p1;

assign mul_ln1352_15_fu_2953_p0 = sext_ln215_15_fu_2825_p1;

assign mul_ln1352_16_fu_2990_p0 = sext_ln215_1_fu_2640_p1;

assign mul_ln1352_17_fu_3003_p0 = sext_ln215_3_fu_2667_p1;

assign mul_ln1352_18_fu_3016_p0 = sext_ln215_5_fu_2694_p1;

assign mul_ln1352_19_fu_3029_p0 = sext_ln215_7_fu_2721_p1;

assign mul_ln1352_1_fu_2671_p0 = sext_ln215_3_fu_2667_p1;

assign mul_ln1352_20_fu_3042_p0 = sext_ln215_9_fu_2748_p1;

assign mul_ln1352_21_fu_3055_p0 = sext_ln215_11_fu_2775_p1;

assign mul_ln1352_22_fu_3064_p0 = sext_ln215_13_fu_2798_p1;

assign mul_ln1352_23_fu_3077_p0 = sext_ln215_15_fu_2825_p1;

assign mul_ln1352_24_fu_3114_p0 = sext_ln215_1_fu_2640_p1;

assign mul_ln1352_25_fu_3127_p0 = sext_ln215_3_fu_2667_p1;

assign mul_ln1352_26_fu_3140_p0 = sext_ln215_5_fu_2694_p1;

assign mul_ln1352_27_fu_3153_p0 = sext_ln215_7_fu_2721_p1;

assign mul_ln1352_28_fu_3166_p0 = sext_ln215_9_fu_2748_p1;

assign mul_ln1352_29_fu_3179_p0 = sext_ln215_11_fu_2775_p1;

assign mul_ln1352_2_fu_2698_p0 = sext_ln215_5_fu_2694_p1;

assign mul_ln1352_30_fu_3188_p0 = sext_ln215_13_fu_2798_p1;

assign mul_ln1352_31_fu_3201_p0 = sext_ln215_15_fu_2825_p1;

assign mul_ln1352_3_fu_2725_p0 = sext_ln215_7_fu_2721_p1;

assign mul_ln1352_4_fu_2752_p0 = sext_ln215_9_fu_2748_p1;

assign mul_ln1352_5_fu_2779_p0 = sext_ln215_11_fu_2775_p1;

assign mul_ln1352_6_fu_2802_p0 = sext_ln215_13_fu_2798_p1;

assign mul_ln1352_7_fu_2829_p0 = sext_ln215_15_fu_2825_p1;

assign mul_ln1352_8_fu_2866_p0 = sext_ln215_1_fu_2640_p1;

assign mul_ln1352_9_fu_2879_p0 = sext_ln215_3_fu_2667_p1;

assign mul_ln1352_fu_2644_p0 = sext_ln215_1_fu_2640_p1;

assign nf_fu_3298_p2 = (nf_assign_fu_708 + 32'd1);

assign out_V_V_TDATA = {{{{add_ln700_83_fu_4825_p2}, {add_ln700_70_fu_4760_p2}}, {add_ln700_57_fu_4695_p2}}, {add_ln700_44_fu_4630_p2}};

assign select_ln271_1_fu_3342_p3 = ((icmp_ln271_reg_5358_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_2_0_fu_440);

assign select_ln271_2_fu_3349_p3 = ((icmp_ln271_reg_5358_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_1_0_fu_436);

assign select_ln271_3_fu_3356_p3 = ((icmp_ln271_reg_5358_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_0_0_fu_432);

assign select_ln271_fu_3335_p3 = ((icmp_ln271_reg_5358_pp0_iter1_reg[0:0] === 1'b1) ? 16'd0 : accu_V_0_3_0_fu_444);

assign select_ln301_fu_3310_p3 = ((icmp_ln301_fu_3304_p2[0:0] === 1'b1) ? 32'd0 : nf_fu_3298_p2);

assign select_ln700_1_fu_4641_p3 = ((xor_ln899_14_fu_4636_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign select_ln700_2_fu_4706_p3 = ((xor_ln899_28_fu_4701_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign select_ln700_3_fu_4771_p3 = ((xor_ln899_42_fu_4766_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign select_ln700_fu_4576_p3 = ((xor_ln899_fu_4571_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign sext_ln170_10_fu_2924_p1 = mul_ln1352_12_fu_2918_p2;

assign sext_ln170_11_fu_2946_p1 = mul_ln1352_14_fu_2940_p2;

assign sext_ln170_12_fu_2996_p1 = mul_ln1352_16_fu_2990_p2;

assign sext_ln170_13_fu_3009_p1 = mul_ln1352_17_fu_3003_p2;

assign sext_ln170_14_fu_3022_p1 = mul_ln1352_18_fu_3016_p2;

assign sext_ln170_15_fu_3035_p1 = mul_ln1352_19_fu_3029_p2;

assign sext_ln170_16_fu_3048_p1 = mul_ln1352_20_fu_3042_p2;

assign sext_ln170_17_fu_3070_p1 = mul_ln1352_22_fu_3064_p2;

assign sext_ln170_18_fu_3120_p1 = mul_ln1352_24_fu_3114_p2;

assign sext_ln170_19_fu_3133_p1 = mul_ln1352_25_fu_3127_p2;

assign sext_ln170_1_fu_2677_p1 = mul_ln1352_1_fu_2671_p2;

assign sext_ln170_20_fu_3146_p1 = mul_ln1352_26_fu_3140_p2;

assign sext_ln170_21_fu_3159_p1 = mul_ln1352_27_fu_3153_p2;

assign sext_ln170_22_fu_3172_p1 = mul_ln1352_28_fu_3166_p2;

assign sext_ln170_23_fu_3194_p1 = mul_ln1352_30_fu_3188_p2;

assign sext_ln170_2_fu_2704_p1 = mul_ln1352_2_fu_2698_p2;

assign sext_ln170_3_fu_2731_p1 = mul_ln1352_3_fu_2725_p2;

assign sext_ln170_4_fu_2758_p1 = mul_ln1352_4_fu_2752_p2;

assign sext_ln170_5_fu_2808_p1 = mul_ln1352_6_fu_2802_p2;

assign sext_ln170_6_fu_2872_p1 = mul_ln1352_8_fu_2866_p2;

assign sext_ln170_7_fu_2885_p1 = mul_ln1352_9_fu_2879_p2;

assign sext_ln170_8_fu_2898_p1 = mul_ln1352_10_fu_2892_p2;

assign sext_ln170_9_fu_2911_p1 = mul_ln1352_11_fu_2905_p2;

assign sext_ln170_fu_2650_p1 = mul_ln1352_fu_2644_p2;

assign sext_ln215_11_fu_2775_p1 = $signed(arg_V_read_assign_5_fu_2762_p4);

assign sext_ln215_13_fu_2798_p1 = $signed(arg_V_read_assign_6_fu_2785_p4);

assign sext_ln215_15_fu_2825_p1 = $signed(arg_V_read_assign_7_fu_2812_p4);

assign sext_ln215_1_fu_2640_p1 = $signed(trunc_ln647_fu_2633_p1);

assign sext_ln215_3_fu_2667_p1 = $signed(arg_V_read_assign_1_fu_2654_p4);

assign sext_ln215_5_fu_2694_p1 = $signed(arg_V_read_assign_2_fu_2681_p4);

assign sext_ln215_7_fu_2721_p1 = $signed(arg_V_read_assign_3_fu_2708_p4);

assign sext_ln215_9_fu_2748_p1 = $signed(arg_V_read_assign_4_fu_2735_p4);

assign sext_ln700_10_fu_3424_p1 = $signed(add_ln700_13_reg_5565);

assign sext_ln700_11_fu_3433_p1 = $signed(add_ln700_14_fu_3427_p2);

assign sext_ln700_12_fu_3443_p1 = mul_ln1352_21_reg_5570;

assign sext_ln700_13_fu_3083_p1 = mul_ln1352_23_fu_3077_p2;

assign sext_ln700_14_fu_3452_p1 = $signed(add_ln700_17_reg_5575);

assign sext_ln700_15_fu_3461_p1 = $signed(add_ln700_19_reg_5580);

assign sext_ln700_16_fu_3464_p1 = $signed(add_ln700_21_reg_5585);

assign sext_ln700_17_fu_3473_p1 = $signed(add_ln700_22_fu_3467_p2);

assign sext_ln700_18_fu_3483_p1 = mul_ln1352_29_reg_5590;

assign sext_ln700_19_fu_3207_p1 = mul_ln1352_31_fu_3201_p2;

assign sext_ln700_1_fu_2835_p1 = mul_ln1352_7_fu_2829_p2;

assign sext_ln700_20_fu_3492_p1 = $signed(add_ln700_25_reg_5595);

assign sext_ln700_21_fu_3501_p1 = $signed(add_ln700_27_reg_5600);

assign sext_ln700_22_fu_3504_p1 = $signed(add_ln700_29_reg_5605);

assign sext_ln700_23_fu_3513_p1 = $signed(add_ln700_30_fu_3507_p2);

assign sext_ln700_2_fu_3372_p1 = $signed(add_ln700_1_reg_5535);

assign sext_ln700_3_fu_3381_p1 = $signed(add_ln700_3_reg_5540);

assign sext_ln700_4_fu_3384_p1 = $signed(add_ln700_5_reg_5545);

assign sext_ln700_5_fu_3393_p1 = $signed(add_ln700_6_fu_3387_p2);

assign sext_ln700_6_fu_3403_p1 = mul_ln1352_13_reg_5550;

assign sext_ln700_7_fu_2959_p1 = mul_ln1352_15_fu_2953_p2;

assign sext_ln700_8_fu_3412_p1 = $signed(add_ln700_9_reg_5555);

assign sext_ln700_9_fu_3421_p1 = $signed(add_ln700_11_reg_5560);

assign sext_ln700_fu_3363_p1 = mul_ln1352_5_reg_5530;

assign sf_fu_2616_p2 = (32'd1 + sf_1_fu_448);

assign threshs_m_thresholds_10_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_11_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_12_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_13_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_14_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_15_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_16_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_17_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_18_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_19_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_1_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_20_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_21_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_22_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_23_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_24_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_25_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_26_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_27_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_28_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_29_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_2_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_30_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_31_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_32_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_33_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_34_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_35_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_36_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_37_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_38_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_39_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_3_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_40_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_41_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_42_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_43_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_44_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_45_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_46_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_47_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_48_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_49_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_4_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_50_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_51_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_52_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_53_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_54_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_55_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_5_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_6_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_7_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_8_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_9_address0 = zext_ln142_fu_3238_p1;

assign threshs_m_thresholds_address0 = zext_ln142_fu_3238_p1;

assign trunc_ln321_fu_1969_p1 = sf_1_fu_448[5:0];

assign trunc_ln647_fu_2633_p1 = ap_phi_reg_pp0_iter1_act_m_val_V_reg_1470[3:0];

assign wgt_M_instance_0_V_fu_2302_p1 = weight_V_V_TDATA[3:0];

assign xor_ln899_10_fu_3942_p2 = (icmp_ln899_10_reg_5940 ^ 1'd1);

assign xor_ln899_11_fu_3951_p2 = (icmp_ln899_11_reg_5945 ^ 1'd1);

assign xor_ln899_12_fu_3960_p2 = (icmp_ln899_12_reg_5950 ^ 1'd1);

assign xor_ln899_13_fu_3969_p2 = (icmp_ln899_13_reg_5955 ^ 1'd1);

assign xor_ln899_14_fu_4636_p2 = (icmp_ln899_14_reg_5960_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_15_fu_4649_p2 = (icmp_ln899_15_reg_5965_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_16_fu_4658_p2 = (icmp_ln899_16_reg_5970_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_17_fu_4052_p2 = (icmp_ln899_17_reg_5975 ^ 1'd1);

assign xor_ln899_18_fu_4061_p2 = (icmp_ln899_18_reg_5980 ^ 1'd1);

assign xor_ln899_19_fu_4070_p2 = (icmp_ln899_19_reg_5985 ^ 1'd1);

assign xor_ln899_1_fu_4584_p2 = (icmp_ln899_1_reg_5895_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_20_fu_4079_p2 = (icmp_ln899_20_reg_5990 ^ 1'd1);

assign xor_ln899_21_fu_4088_p2 = (icmp_ln899_21_reg_5995 ^ 1'd1);

assign xor_ln899_22_fu_4097_p2 = (icmp_ln899_22_reg_6000 ^ 1'd1);

assign xor_ln899_23_fu_4106_p2 = (icmp_ln899_23_reg_6005 ^ 1'd1);

assign xor_ln899_24_fu_4115_p2 = (icmp_ln899_24_reg_6010 ^ 1'd1);

assign xor_ln899_25_fu_4124_p2 = (icmp_ln899_25_reg_6015 ^ 1'd1);

assign xor_ln899_26_fu_4133_p2 = (icmp_ln899_26_reg_6020 ^ 1'd1);

assign xor_ln899_27_fu_4142_p2 = (icmp_ln899_27_reg_6025 ^ 1'd1);

assign xor_ln899_28_fu_4701_p2 = (icmp_ln899_28_reg_6030_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_29_fu_4714_p2 = (icmp_ln899_29_reg_6035_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_2_fu_4593_p2 = (icmp_ln899_2_reg_5900_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_30_fu_4723_p2 = (icmp_ln899_30_reg_6040_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_31_fu_4225_p2 = (icmp_ln899_31_reg_6045 ^ 1'd1);

assign xor_ln899_32_fu_4234_p2 = (icmp_ln899_32_reg_6050 ^ 1'd1);

assign xor_ln899_33_fu_4243_p2 = (icmp_ln899_33_reg_6055 ^ 1'd1);

assign xor_ln899_34_fu_4252_p2 = (icmp_ln899_34_reg_6060 ^ 1'd1);

assign xor_ln899_35_fu_4261_p2 = (icmp_ln899_35_reg_6065 ^ 1'd1);

assign xor_ln899_36_fu_4270_p2 = (icmp_ln899_36_reg_6070 ^ 1'd1);

assign xor_ln899_37_fu_4279_p2 = (icmp_ln899_37_reg_6075 ^ 1'd1);

assign xor_ln899_38_fu_4288_p2 = (icmp_ln899_38_reg_6080 ^ 1'd1);

assign xor_ln899_39_fu_4297_p2 = (icmp_ln899_39_reg_6085 ^ 1'd1);

assign xor_ln899_3_fu_3879_p2 = (icmp_ln899_3_reg_5905 ^ 1'd1);

assign xor_ln899_40_fu_4306_p2 = (icmp_ln899_40_reg_6090 ^ 1'd1);

assign xor_ln899_41_fu_4315_p2 = (icmp_ln899_41_reg_6095 ^ 1'd1);

assign xor_ln899_42_fu_4766_p2 = (icmp_ln899_42_reg_6100_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_43_fu_4779_p2 = (icmp_ln899_43_reg_6105_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_44_fu_4788_p2 = (icmp_ln899_44_reg_6110_pp0_iter3_reg ^ 1'd1);

assign xor_ln899_45_fu_4398_p2 = (icmp_ln899_45_reg_6115 ^ 1'd1);

assign xor_ln899_46_fu_4407_p2 = (icmp_ln899_46_reg_6120 ^ 1'd1);

assign xor_ln899_47_fu_4416_p2 = (icmp_ln899_47_reg_6125 ^ 1'd1);

assign xor_ln899_48_fu_4425_p2 = (icmp_ln899_48_reg_6130 ^ 1'd1);

assign xor_ln899_49_fu_4434_p2 = (icmp_ln899_49_reg_6135 ^ 1'd1);

assign xor_ln899_4_fu_3888_p2 = (icmp_ln899_4_reg_5910 ^ 1'd1);

assign xor_ln899_50_fu_4443_p2 = (icmp_ln899_50_reg_6140 ^ 1'd1);

assign xor_ln899_51_fu_4452_p2 = (icmp_ln899_51_reg_6145 ^ 1'd1);

assign xor_ln899_52_fu_4461_p2 = (icmp_ln899_52_reg_6150 ^ 1'd1);

assign xor_ln899_53_fu_4470_p2 = (icmp_ln899_53_reg_6155 ^ 1'd1);

assign xor_ln899_54_fu_4479_p2 = (icmp_ln899_54_reg_6160 ^ 1'd1);

assign xor_ln899_55_fu_4488_p2 = (icmp_ln899_55_reg_6165 ^ 1'd1);

assign xor_ln899_5_fu_3897_p2 = (icmp_ln899_5_reg_5915 ^ 1'd1);

assign xor_ln899_6_fu_3906_p2 = (icmp_ln899_6_reg_5920 ^ 1'd1);

assign xor_ln899_7_fu_3915_p2 = (icmp_ln899_7_reg_5925 ^ 1'd1);

assign xor_ln899_8_fu_3924_p2 = (icmp_ln899_8_reg_5930 ^ 1'd1);

assign xor_ln899_9_fu_3933_p2 = (icmp_ln899_9_reg_5935 ^ 1'd1);

assign xor_ln899_fu_4571_p2 = (icmp_ln899_reg_5890_pp0_iter3_reg ^ 1'd1);

assign zext_ln142_10_fu_3947_p1 = xor_ln899_10_fu_3942_p2;

assign zext_ln142_11_fu_3956_p1 = xor_ln899_11_fu_3951_p2;

assign zext_ln142_12_fu_3965_p1 = xor_ln899_12_fu_3960_p2;

assign zext_ln142_13_fu_4654_p1 = xor_ln899_15_fu_4649_p2;

assign zext_ln142_14_fu_4663_p1 = xor_ln899_16_fu_4658_p2;

assign zext_ln142_15_fu_4057_p1 = xor_ln899_17_fu_4052_p2;

assign zext_ln142_16_fu_4066_p1 = xor_ln899_18_fu_4061_p2;

assign zext_ln142_17_fu_4075_p1 = xor_ln899_19_fu_4070_p2;

assign zext_ln142_18_fu_4084_p1 = xor_ln899_20_fu_4079_p2;

assign zext_ln142_19_fu_4093_p1 = xor_ln899_21_fu_4088_p2;

assign zext_ln142_1_fu_4589_p1 = xor_ln899_1_fu_4584_p2;

assign zext_ln142_20_fu_4102_p1 = xor_ln899_22_fu_4097_p2;

assign zext_ln142_21_fu_4111_p1 = xor_ln899_23_fu_4106_p2;

assign zext_ln142_22_fu_4120_p1 = xor_ln899_24_fu_4115_p2;

assign zext_ln142_23_fu_4129_p1 = xor_ln899_25_fu_4124_p2;

assign zext_ln142_24_fu_4138_p1 = xor_ln899_26_fu_4133_p2;

assign zext_ln142_25_fu_4719_p1 = xor_ln899_29_fu_4714_p2;

assign zext_ln142_26_fu_4728_p1 = xor_ln899_30_fu_4723_p2;

assign zext_ln142_27_fu_4230_p1 = xor_ln899_31_fu_4225_p2;

assign zext_ln142_28_fu_4239_p1 = xor_ln899_32_fu_4234_p2;

assign zext_ln142_29_fu_4248_p1 = xor_ln899_33_fu_4243_p2;

assign zext_ln142_2_fu_4598_p1 = xor_ln899_2_fu_4593_p2;

assign zext_ln142_30_fu_4257_p1 = xor_ln899_34_fu_4252_p2;

assign zext_ln142_31_fu_4266_p1 = xor_ln899_35_fu_4261_p2;

assign zext_ln142_32_fu_4275_p1 = xor_ln899_36_fu_4270_p2;

assign zext_ln142_33_fu_4284_p1 = xor_ln899_37_fu_4279_p2;

assign zext_ln142_34_fu_4293_p1 = xor_ln899_38_fu_4288_p2;

assign zext_ln142_35_fu_4302_p1 = xor_ln899_39_fu_4297_p2;

assign zext_ln142_36_fu_4311_p1 = xor_ln899_40_fu_4306_p2;

assign zext_ln142_37_fu_4784_p1 = xor_ln899_43_fu_4779_p2;

assign zext_ln142_38_fu_4793_p1 = xor_ln899_44_fu_4788_p2;

assign zext_ln142_39_fu_4403_p1 = xor_ln899_45_fu_4398_p2;

assign zext_ln142_3_fu_3884_p1 = xor_ln899_3_fu_3879_p2;

assign zext_ln142_40_fu_4412_p1 = xor_ln899_46_fu_4407_p2;

assign zext_ln142_41_fu_4421_p1 = xor_ln899_47_fu_4416_p2;

assign zext_ln142_42_fu_4430_p1 = xor_ln899_48_fu_4425_p2;

assign zext_ln142_43_fu_4439_p1 = xor_ln899_49_fu_4434_p2;

assign zext_ln142_44_fu_4448_p1 = xor_ln899_50_fu_4443_p2;

assign zext_ln142_45_fu_4457_p1 = xor_ln899_51_fu_4452_p2;

assign zext_ln142_46_fu_4466_p1 = xor_ln899_52_fu_4461_p2;

assign zext_ln142_47_fu_4475_p1 = xor_ln899_53_fu_4470_p2;

assign zext_ln142_48_fu_4484_p1 = xor_ln899_54_fu_4479_p2;

assign zext_ln142_4_fu_3893_p1 = xor_ln899_4_fu_3888_p2;

assign zext_ln142_5_fu_3902_p1 = xor_ln899_5_fu_3897_p2;

assign zext_ln142_6_fu_3911_p1 = xor_ln899_6_fu_3906_p2;

assign zext_ln142_7_fu_3920_p1 = xor_ln899_7_fu_3915_p2;

assign zext_ln142_8_fu_3929_p1 = xor_ln899_8_fu_3924_p2;

assign zext_ln142_9_fu_3938_p1 = xor_ln899_9_fu_3933_p2;

assign zext_ln142_fu_3238_p1 = nf_assign_fu_708;

assign zext_ln700_10_fu_4673_p1 = add_ln700_45_fu_4667_p2;

assign zext_ln700_11_fu_4157_p1 = add_ln700_47_fu_4151_p2;

assign zext_ln700_12_fu_4167_p1 = add_ln700_48_fu_4161_p2;

assign zext_ln700_13_fu_4683_p1 = add_ln700_49_reg_6180;

assign zext_ln700_14_fu_4189_p1 = add_ln700_52_fu_4183_p2;

assign zext_ln700_15_fu_4199_p1 = add_ln700_53_fu_4193_p2;

assign zext_ln700_16_fu_4209_p1 = add_ln700_54_fu_4203_p2;

assign zext_ln700_17_fu_4692_p1 = add_ln700_56_reg_6185;

assign zext_ln700_18_fu_4320_p1 = xor_ln899_41_fu_4315_p2;

assign zext_ln700_19_fu_4738_p1 = add_ln700_58_fu_4732_p2;

assign zext_ln700_1_fu_4608_p1 = add_ln700_32_fu_4602_p2;

assign zext_ln700_20_fu_4330_p1 = add_ln700_60_fu_4324_p2;

assign zext_ln700_21_fu_4340_p1 = add_ln700_61_fu_4334_p2;

assign zext_ln700_22_fu_4748_p1 = add_ln700_62_reg_6190;

assign zext_ln700_23_fu_4362_p1 = add_ln700_65_fu_4356_p2;

assign zext_ln700_24_fu_4372_p1 = add_ln700_66_fu_4366_p2;

assign zext_ln700_25_fu_4382_p1 = add_ln700_67_fu_4376_p2;

assign zext_ln700_26_fu_4757_p1 = add_ln700_69_reg_6195;

assign zext_ln700_27_fu_4493_p1 = xor_ln899_55_fu_4488_p2;

assign zext_ln700_28_fu_4803_p1 = add_ln700_71_fu_4797_p2;

assign zext_ln700_29_fu_4503_p1 = add_ln700_73_fu_4497_p2;

assign zext_ln700_2_fu_3984_p1 = add_ln700_34_fu_3978_p2;

assign zext_ln700_30_fu_4513_p1 = add_ln700_74_fu_4507_p2;

assign zext_ln700_31_fu_4813_p1 = add_ln700_75_reg_6200;

assign zext_ln700_32_fu_4535_p1 = add_ln700_78_fu_4529_p2;

assign zext_ln700_33_fu_4545_p1 = add_ln700_79_fu_4539_p2;

assign zext_ln700_34_fu_4555_p1 = add_ln700_80_fu_4549_p2;

assign zext_ln700_35_fu_4822_p1 = add_ln700_82_reg_6205;

assign zext_ln700_3_fu_3994_p1 = add_ln700_35_fu_3988_p2;

assign zext_ln700_4_fu_4618_p1 = add_ln700_36_reg_6170;

assign zext_ln700_5_fu_4016_p1 = add_ln700_39_fu_4010_p2;

assign zext_ln700_6_fu_4026_p1 = add_ln700_40_fu_4020_p2;

assign zext_ln700_7_fu_4036_p1 = add_ln700_41_fu_4030_p2;

assign zext_ln700_8_fu_4627_p1 = add_ln700_43_reg_6175;

assign zext_ln700_9_fu_4147_p1 = xor_ln899_27_fu_4142_p2;

assign zext_ln700_fu_3974_p1 = xor_ln899_13_fu_3969_p2;

endmodule //StreamingFCLayer_Batch_4_Matrix_Vector_Activa
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_StreamingFCLayer_Batch_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingFCLayer_Batch_1_StreamingFCLayer_Batch_1,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=8.042250,HLS_SYN_LAT=36871,HLS_SYN_TPT=none,HLS_SYN_MEM=56,HLS_SYN_DSP=0,HLS_SYN_FF=9651,HLS_SYN_LUT=5149,HLS_VERSION=2020_1_1}" *)

module StreamingFCLayer_Batch_1_StreamingFCLayer_Batch_1 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        weights_V_V_TDATA,
        weights_V_V_TVALID,
        weights_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
input  [63:0] weights_V_V_TDATA;
input   weights_V_V_TVALID;
output   weights_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;
reg weights_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_Matrix_Vector_Activa_fu_140_ap_start;
wire    grp_Matrix_Vector_Activa_fu_140_ap_done;
wire    grp_Matrix_Vector_Activa_fu_140_ap_idle;
wire    grp_Matrix_Vector_Activa_fu_140_ap_ready;
wire    grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY;
wire   [15:0] grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA;
wire    grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID;
wire    grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY;
wire    grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY;
reg    grp_Matrix_Vector_Activa_fu_140_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [15:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    regslice_both_weights_V_V_U_apdone_blk;
wire   [63:0] weights_V_V_TDATA_int;
wire    weights_V_V_TVALID_int;
reg    weights_V_V_TREADY_int;
wire    regslice_both_weights_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_Matrix_Vector_Activa_fu_140_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingFCLayer_Batch_1_Matrix_Vector_Activa grp_Matrix_Vector_Activa_fu_140(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_Matrix_Vector_Activa_fu_140_ap_start),
    .ap_done(grp_Matrix_Vector_Activa_fu_140_ap_done),
    .ap_idle(grp_Matrix_Vector_Activa_fu_140_ap_idle),
    .ap_ready(grp_Matrix_Vector_Activa_fu_140_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY),
    .out_V_V_TDATA(grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA),
    .out_V_V_TVALID(grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID),
    .out_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY),
    .weight_V_V_TDATA(weights_V_V_TDATA_int),
    .weight_V_V_TVALID(weights_V_V_TVALID_int),
    .weight_V_V_TREADY(grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 64 ))
regslice_both_weights_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(weights_V_V_TDATA),
    .vld_in(weights_V_V_TVALID),
    .ack_in(regslice_both_weights_V_V_U_ack_in),
    .data_out(weights_V_V_TDATA_int),
    .vld_out(weights_V_V_TVALID_int),
    .ack_out(weights_V_V_TREADY_int),
    .apdone_blk(regslice_both_weights_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_Matrix_Vector_Activa_fu_140_out_V_V_TDATA),
    .vld_in(grp_Matrix_Vector_Activa_fu_140_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b1;
        end else if ((grp_Matrix_Vector_Activa_fu_140_ap_ready == 1'b1)) begin
            grp_Matrix_Vector_Activa_fu_140_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_140_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    if (((regslice_both_weights_V_V_U_ack_in == 1'b1) & (weights_V_V_TVALID == 1'b1))) begin
        weights_V_V_TREADY = 1'b1;
    end else begin
        weights_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        weights_V_V_TREADY_int = grp_Matrix_Vector_Activa_fu_140_weight_V_V_TREADY;
    end else begin
        weights_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_Matrix_Vector_Activa_fu_140_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_Matrix_Vector_Activa_fu_140_ap_start = grp_Matrix_Vector_Activa_fu_140_ap_start_reg;

assign grp_Matrix_Vector_Activa_fu_140_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingFCLayer_Batch_1_StreamingFCLayer_Batch_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcclv.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcclv_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcclv_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcclv(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcclv_rom Thresholding_Batch_0_Thresholding_Batcclv_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actyd2.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actyd2_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actyd2_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actyd2(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actyd2_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actyd2_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcocq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_Batcocq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcocq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_Batcocq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_Batcocq_rom Thresholding_Batch_2_Thresholding_Batcocq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/synth/finn_design.v

//Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
//--------------------------------------------------------------------------------
//Tool Version: Vivado v.2020.1.1 (lin64) Build 2960000 Wed Aug  5 22:57:21 MDT 2020
//Date        : Sat Jan 30 13:23:55 2021
//Host        : finn_dev_grgov running 64-bit unknown
//Command     : generate_target finn_design.bd
//Design      : finn_design
//Purpose     : IP block netlist
//--------------------------------------------------------------------------------
`timescale 1 ps / 1 ps

module StreamingFCLayer_Batch_0_imp_5FXKV0
   (ap_clk,
    ap_rst_n,
    in0_V_V_tdata,
    in0_V_V_tready,
    in0_V_V_tvalid,
    out_V_V_tdata,
    out_V_V_tready,
    out_V_V_tvalid);
  input ap_clk;
  input ap_rst_n;
  input [7:0]in0_V_V_tdata;
  output in0_V_V_tready;
  input in0_V_V_tvalid;
  output [95:0]out_V_V_tdata;
  input out_V_V_tready;
  output out_V_V_tvalid;

  wire [95:0]StreamingFCLayer_Batch_0_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_0_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_0_out_V_V_TVALID;
  wire [31:0]StreamingFCLayer_Batch_0_wstrm_m_axis_0_TDATA;
  wire StreamingFCLayer_Batch_0_wstrm_m_axis_0_TREADY;
  wire StreamingFCLayer_Batch_0_wstrm_m_axis_0_TVALID;
  wire ap_clk_1;
  wire ap_rst_n_1;
  wire [7:0]in0_V_V_1_TDATA;
  wire in0_V_V_1_TREADY;
  wire in0_V_V_1_TVALID;

  assign StreamingFCLayer_Batch_0_out_V_V_TREADY = out_V_V_tready;
  assign ap_clk_1 = ap_clk;
  assign ap_rst_n_1 = ap_rst_n;
  assign in0_V_V_1_TDATA = in0_V_V_tdata[7:0];
  assign in0_V_V_1_TVALID = in0_V_V_tvalid;
  assign in0_V_V_tready = in0_V_V_1_TREADY;
  assign out_V_V_tdata[95:0] = StreamingFCLayer_Batch_0_out_V_V_TDATA;
  assign out_V_V_tvalid = StreamingFCLayer_Batch_0_out_V_V_TVALID;
  finn_design_StreamingFCLayer_Batch_0_0 StreamingFCLayer_Batch_0
       (.ap_clk(ap_clk_1),
        .ap_rst_n(ap_rst_n_1),
        .in0_V_V_TDATA(in0_V_V_1_TDATA),
        .in0_V_V_TREADY(in0_V_V_1_TREADY),
        .in0_V_V_TVALID(in0_V_V_1_TVALID),
        .out_V_V_TDATA(StreamingFCLayer_Batch_0_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFCLayer_Batch_0_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFCLayer_Batch_0_out_V_V_TVALID),
        .weights_V_V_TDATA(StreamingFCLayer_Batch_0_wstrm_m_axis_0_TDATA),
        .weights_V_V_TREADY(StreamingFCLayer_Batch_0_wstrm_m_axis_0_TREADY),
        .weights_V_V_TVALID(StreamingFCLayer_Batch_0_wstrm_m_axis_0_TVALID));
  finn_design_StreamingFCLayer_Batch_0_wstrm_0 StreamingFCLayer_Batch_0_wstrm
       (.aclk(ap_clk_1),
        .araddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .aresetn(ap_rst_n_1),
        .arprot({1'b0,1'b0,1'b0}),
        .arvalid(1'b0),
        .awaddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .awprot({1'b0,1'b0,1'b0}),
        .awvalid(1'b0),
        .bready(1'b0),
        .m_axis_0_tdata(StreamingFCLayer_Batch_0_wstrm_m_axis_0_TDATA),
        .m_axis_0_tready(StreamingFCLayer_Batch_0_wstrm_m_axis_0_TREADY),
        .m_axis_0_tvalid(StreamingFCLayer_Batch_0_wstrm_m_axis_0_TVALID),
        .rready(1'b0),
        .wdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .wstrb({1'b1,1'b1,1'b1,1'b1}),
        .wvalid(1'b0));
endmodule

module StreamingFCLayer_Batch_1_imp_11SOJ3N
   (ap_clk,
    ap_rst_n,
    in0_V_V_tdata,
    in0_V_V_tready,
    in0_V_V_tvalid,
    out_V_V_tdata,
    out_V_V_tready,
    out_V_V_tvalid);
  input ap_clk;
  input ap_rst_n;
  input [15:0]in0_V_V_tdata;
  output in0_V_V_tready;
  input in0_V_V_tvalid;
  output [15:0]out_V_V_tdata;
  input out_V_V_tready;
  output out_V_V_tvalid;

  wire [15:0]StreamingFCLayer_Batch_1_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_1_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_1_out_V_V_TVALID;
  wire [63:0]StreamingFCLayer_Batch_1_wstrm_m_axis_0_TDATA;
  wire StreamingFCLayer_Batch_1_wstrm_m_axis_0_TREADY;
  wire StreamingFCLayer_Batch_1_wstrm_m_axis_0_TVALID;
  wire ap_clk_1;
  wire ap_rst_n_1;
  wire [15:0]in0_V_V_1_TDATA;
  wire in0_V_V_1_TREADY;
  wire in0_V_V_1_TVALID;

  assign StreamingFCLayer_Batch_1_out_V_V_TREADY = out_V_V_tready;
  assign ap_clk_1 = ap_clk;
  assign ap_rst_n_1 = ap_rst_n;
  assign in0_V_V_1_TDATA = in0_V_V_tdata[15:0];
  assign in0_V_V_1_TVALID = in0_V_V_tvalid;
  assign in0_V_V_tready = in0_V_V_1_TREADY;
  assign out_V_V_tdata[15:0] = StreamingFCLayer_Batch_1_out_V_V_TDATA;
  assign out_V_V_tvalid = StreamingFCLayer_Batch_1_out_V_V_TVALID;
  finn_design_StreamingFCLayer_Batch_1_0 StreamingFCLayer_Batch_1
       (.ap_clk(ap_clk_1),
        .ap_rst_n(ap_rst_n_1),
        .in0_V_V_TDATA(in0_V_V_1_TDATA),
        .in0_V_V_TREADY(in0_V_V_1_TREADY),
        .in0_V_V_TVALID(in0_V_V_1_TVALID),
        .out_V_V_TDATA(StreamingFCLayer_Batch_1_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFCLayer_Batch_1_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFCLayer_Batch_1_out_V_V_TVALID),
        .weights_V_V_TDATA(StreamingFCLayer_Batch_1_wstrm_m_axis_0_TDATA),
        .weights_V_V_TREADY(StreamingFCLayer_Batch_1_wstrm_m_axis_0_TREADY),
        .weights_V_V_TVALID(StreamingFCLayer_Batch_1_wstrm_m_axis_0_TVALID));
  finn_design_StreamingFCLayer_Batch_1_wstrm_0 StreamingFCLayer_Batch_1_wstrm
       (.aclk(ap_clk_1),
        .araddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .aresetn(ap_rst_n_1),
        .arprot({1'b0,1'b0,1'b0}),
        .arvalid(1'b0),
        .awaddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .awprot({1'b0,1'b0,1'b0}),
        .awvalid(1'b0),
        .bready(1'b0),
        .m_axis_0_tdata(StreamingFCLayer_Batch_1_wstrm_m_axis_0_TDATA),
        .m_axis_0_tready(StreamingFCLayer_Batch_1_wstrm_m_axis_0_TREADY),
        .m_axis_0_tvalid(StreamingFCLayer_Batch_1_wstrm_m_axis_0_TVALID),
        .rready(1'b0),
        .wdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .wstrb({1'b1,1'b1,1'b1,1'b1}),
        .wvalid(1'b0));
endmodule

module StreamingFCLayer_Batch_2_imp_1YXLQV7
   (ap_clk,
    ap_rst_n,
    in0_V_V_tdata,
    in0_V_V_tready,
    in0_V_V_tvalid,
    out_V_V_tdata,
    out_V_V_tready,
    out_V_V_tvalid);
  input ap_clk;
  input ap_rst_n;
  input [31:0]in0_V_V_tdata;
  output in0_V_V_tready;
  input in0_V_V_tvalid;
  output [15:0]out_V_V_tdata;
  input out_V_V_tready;
  output out_V_V_tvalid;

  wire [15:0]StreamingFCLayer_Batch_2_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_2_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_2_out_V_V_TVALID;
  wire [127:0]StreamingFCLayer_Batch_2_wstrm_m_axis_0_TDATA;
  wire StreamingFCLayer_Batch_2_wstrm_m_axis_0_TREADY;
  wire StreamingFCLayer_Batch_2_wstrm_m_axis_0_TVALID;
  wire ap_clk_1;
  wire ap_rst_n_1;
  wire [31:0]in0_V_V_1_TDATA;
  wire in0_V_V_1_TREADY;
  wire in0_V_V_1_TVALID;

  assign StreamingFCLayer_Batch_2_out_V_V_TREADY = out_V_V_tready;
  assign ap_clk_1 = ap_clk;
  assign ap_rst_n_1 = ap_rst_n;
  assign in0_V_V_1_TDATA = in0_V_V_tdata[31:0];
  assign in0_V_V_1_TVALID = in0_V_V_tvalid;
  assign in0_V_V_tready = in0_V_V_1_TREADY;
  assign out_V_V_tdata[15:0] = StreamingFCLayer_Batch_2_out_V_V_TDATA;
  assign out_V_V_tvalid = StreamingFCLayer_Batch_2_out_V_V_TVALID;
  finn_design_StreamingFCLayer_Batch_2_0 StreamingFCLayer_Batch_2
       (.ap_clk(ap_clk_1),
        .ap_rst_n(ap_rst_n_1),
        .in0_V_V_TDATA(in0_V_V_1_TDATA),
        .in0_V_V_TREADY(in0_V_V_1_TREADY),
        .in0_V_V_TVALID(in0_V_V_1_TVALID),
        .out_V_V_TDATA(StreamingFCLayer_Batch_2_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFCLayer_Batch_2_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFCLayer_Batch_2_out_V_V_TVALID),
        .weights_V_V_TDATA(StreamingFCLayer_Batch_2_wstrm_m_axis_0_TDATA),
        .weights_V_V_TREADY(StreamingFCLayer_Batch_2_wstrm_m_axis_0_TREADY),
        .weights_V_V_TVALID(StreamingFCLayer_Batch_2_wstrm_m_axis_0_TVALID));
  finn_design_StreamingFCLayer_Batch_2_wstrm_0 StreamingFCLayer_Batch_2_wstrm
       (.aclk(ap_clk_1),
        .araddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .aresetn(ap_rst_n_1),
        .arprot({1'b0,1'b0,1'b0}),
        .arvalid(1'b0),
        .awaddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .awprot({1'b0,1'b0,1'b0}),
        .awvalid(1'b0),
        .bready(1'b0),
        .m_axis_0_tdata(StreamingFCLayer_Batch_2_wstrm_m_axis_0_TDATA),
        .m_axis_0_tready(StreamingFCLayer_Batch_2_wstrm_m_axis_0_TREADY),
        .m_axis_0_tvalid(StreamingFCLayer_Batch_2_wstrm_m_axis_0_TVALID),
        .rready(1'b0),
        .wdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .wstrb({1'b1,1'b1,1'b1,1'b1}),
        .wvalid(1'b0));
endmodule

module StreamingFCLayer_Batch_3_imp_RR03E4
   (ap_clk,
    ap_rst_n,
    in0_V_V_tdata,
    in0_V_V_tready,
    in0_V_V_tvalid,
    out_V_V_tdata,
    out_V_V_tready,
    out_V_V_tvalid);
  input ap_clk;
  input ap_rst_n;
  input [23:0]in0_V_V_tdata;
  output in0_V_V_tready;
  input in0_V_V_tvalid;
  output [15:0]out_V_V_tdata;
  input out_V_V_tready;
  output out_V_V_tvalid;

  wire [15:0]StreamingFCLayer_Batch_3_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_3_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_3_out_V_V_TVALID;
  wire [47:0]StreamingFCLayer_Batch_3_wstrm_m_axis_0_TDATA;
  wire StreamingFCLayer_Batch_3_wstrm_m_axis_0_TREADY;
  wire StreamingFCLayer_Batch_3_wstrm_m_axis_0_TVALID;
  wire ap_clk_1;
  wire ap_rst_n_1;
  wire [23:0]in0_V_V_1_TDATA;
  wire in0_V_V_1_TREADY;
  wire in0_V_V_1_TVALID;

  assign StreamingFCLayer_Batch_3_out_V_V_TREADY = out_V_V_tready;
  assign ap_clk_1 = ap_clk;
  assign ap_rst_n_1 = ap_rst_n;
  assign in0_V_V_1_TDATA = in0_V_V_tdata[23:0];
  assign in0_V_V_1_TVALID = in0_V_V_tvalid;
  assign in0_V_V_tready = in0_V_V_1_TREADY;
  assign out_V_V_tdata[15:0] = StreamingFCLayer_Batch_3_out_V_V_TDATA;
  assign out_V_V_tvalid = StreamingFCLayer_Batch_3_out_V_V_TVALID;
  finn_design_StreamingFCLayer_Batch_3_0 StreamingFCLayer_Batch_3
       (.ap_clk(ap_clk_1),
        .ap_rst_n(ap_rst_n_1),
        .in0_V_V_TDATA(in0_V_V_1_TDATA),
        .in0_V_V_TREADY(in0_V_V_1_TREADY),
        .in0_V_V_TVALID(in0_V_V_1_TVALID),
        .out_V_V_TDATA(StreamingFCLayer_Batch_3_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFCLayer_Batch_3_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFCLayer_Batch_3_out_V_V_TVALID),
        .weights_V_V_TDATA(StreamingFCLayer_Batch_3_wstrm_m_axis_0_TDATA),
        .weights_V_V_TREADY(StreamingFCLayer_Batch_3_wstrm_m_axis_0_TREADY),
        .weights_V_V_TVALID(StreamingFCLayer_Batch_3_wstrm_m_axis_0_TVALID));
  finn_design_StreamingFCLayer_Batch_3_wstrm_0 StreamingFCLayer_Batch_3_wstrm
       (.aclk(ap_clk_1),
        .araddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .aresetn(ap_rst_n_1),
        .arprot({1'b0,1'b0,1'b0}),
        .arvalid(1'b0),
        .awaddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .awprot({1'b0,1'b0,1'b0}),
        .awvalid(1'b0),
        .bready(1'b0),
        .m_axis_0_tdata(StreamingFCLayer_Batch_3_wstrm_m_axis_0_TDATA),
        .m_axis_0_tready(StreamingFCLayer_Batch_3_wstrm_m_axis_0_TREADY),
        .m_axis_0_tvalid(StreamingFCLayer_Batch_3_wstrm_m_axis_0_TVALID),
        .rready(1'b0),
        .wdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .wstrb({1'b1,1'b1,1'b1,1'b1}),
        .wvalid(1'b0));
endmodule

module StreamingFCLayer_Batch_4_imp_4LW78J
   (ap_clk,
    ap_rst_n,
    in0_V_V_tdata,
    in0_V_V_tready,
    in0_V_V_tvalid,
    out_V_V_tdata,
    out_V_V_tready,
    out_V_V_tvalid);
  input ap_clk;
  input ap_rst_n;
  input [31:0]in0_V_V_tdata;
  output in0_V_V_tready;
  input in0_V_V_tvalid;
  output [15:0]out_V_V_tdata;
  input out_V_V_tready;
  output out_V_V_tvalid;

  wire [15:0]StreamingFCLayer_Batch_4_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_4_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_4_out_V_V_TVALID;
  wire [127:0]StreamingFCLayer_Batch_4_wstrm_m_axis_0_TDATA;
  wire StreamingFCLayer_Batch_4_wstrm_m_axis_0_TREADY;
  wire StreamingFCLayer_Batch_4_wstrm_m_axis_0_TVALID;
  wire ap_clk_1;
  wire ap_rst_n_1;
  wire [31:0]in0_V_V_1_TDATA;
  wire in0_V_V_1_TREADY;
  wire in0_V_V_1_TVALID;

  assign StreamingFCLayer_Batch_4_out_V_V_TREADY = out_V_V_tready;
  assign ap_clk_1 = ap_clk;
  assign ap_rst_n_1 = ap_rst_n;
  assign in0_V_V_1_TDATA = in0_V_V_tdata[31:0];
  assign in0_V_V_1_TVALID = in0_V_V_tvalid;
  assign in0_V_V_tready = in0_V_V_1_TREADY;
  assign out_V_V_tdata[15:0] = StreamingFCLayer_Batch_4_out_V_V_TDATA;
  assign out_V_V_tvalid = StreamingFCLayer_Batch_4_out_V_V_TVALID;
  finn_design_StreamingFCLayer_Batch_4_0 StreamingFCLayer_Batch_4
       (.ap_clk(ap_clk_1),
        .ap_rst_n(ap_rst_n_1),
        .in0_V_V_TDATA(in0_V_V_1_TDATA),
        .in0_V_V_TREADY(in0_V_V_1_TREADY),
        .in0_V_V_TVALID(in0_V_V_1_TVALID),
        .out_V_V_TDATA(StreamingFCLayer_Batch_4_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFCLayer_Batch_4_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFCLayer_Batch_4_out_V_V_TVALID),
        .weights_V_V_TDATA(StreamingFCLayer_Batch_4_wstrm_m_axis_0_TDATA),
        .weights_V_V_TREADY(StreamingFCLayer_Batch_4_wstrm_m_axis_0_TREADY),
        .weights_V_V_TVALID(StreamingFCLayer_Batch_4_wstrm_m_axis_0_TVALID));
  finn_design_StreamingFCLayer_Batch_4_wstrm_0 StreamingFCLayer_Batch_4_wstrm
       (.aclk(ap_clk_1),
        .araddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .aresetn(ap_rst_n_1),
        .arprot({1'b0,1'b0,1'b0}),
        .arvalid(1'b0),
        .awaddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .awprot({1'b0,1'b0,1'b0}),
        .awvalid(1'b0),
        .bready(1'b0),
        .m_axis_0_tdata(StreamingFCLayer_Batch_4_wstrm_m_axis_0_TDATA),
        .m_axis_0_tready(StreamingFCLayer_Batch_4_wstrm_m_axis_0_TREADY),
        .m_axis_0_tvalid(StreamingFCLayer_Batch_4_wstrm_m_axis_0_TVALID),
        .rready(1'b0),
        .wdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .wstrb({1'b1,1'b1,1'b1,1'b1}),
        .wvalid(1'b0));
endmodule

module StreamingFCLayer_Batch_5_imp_12MW1JG
   (ap_clk,
    ap_rst_n,
    in0_V_V_tdata,
    in0_V_V_tready,
    in0_V_V_tvalid,
    out_V_V_tdata,
    out_V_V_tready,
    out_V_V_tvalid);
  input ap_clk;
  input ap_rst_n;
  input [31:0]in0_V_V_tdata;
  output in0_V_V_tready;
  input in0_V_V_tvalid;
  output [15:0]out_V_V_tdata;
  input out_V_V_tready;
  output out_V_V_tvalid;

  wire [15:0]StreamingFCLayer_Batch_5_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_5_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_5_out_V_V_TVALID;
  wire [31:0]StreamingFCLayer_Batch_5_wstrm_m_axis_0_TDATA;
  wire StreamingFCLayer_Batch_5_wstrm_m_axis_0_TREADY;
  wire StreamingFCLayer_Batch_5_wstrm_m_axis_0_TVALID;
  wire ap_clk_1;
  wire ap_rst_n_1;
  wire [31:0]in0_V_V_1_TDATA;
  wire in0_V_V_1_TREADY;
  wire in0_V_V_1_TVALID;

  assign StreamingFCLayer_Batch_5_out_V_V_TREADY = out_V_V_tready;
  assign ap_clk_1 = ap_clk;
  assign ap_rst_n_1 = ap_rst_n;
  assign in0_V_V_1_TDATA = in0_V_V_tdata[31:0];
  assign in0_V_V_1_TVALID = in0_V_V_tvalid;
  assign in0_V_V_tready = in0_V_V_1_TREADY;
  assign out_V_V_tdata[15:0] = StreamingFCLayer_Batch_5_out_V_V_TDATA;
  assign out_V_V_tvalid = StreamingFCLayer_Batch_5_out_V_V_TVALID;
  finn_design_StreamingFCLayer_Batch_5_0 StreamingFCLayer_Batch_5
       (.ap_clk(ap_clk_1),
        .ap_rst_n(ap_rst_n_1),
        .in0_V_V_TDATA(in0_V_V_1_TDATA),
        .in0_V_V_TREADY(in0_V_V_1_TREADY),
        .in0_V_V_TVALID(in0_V_V_1_TVALID),
        .out_V_V_TDATA(StreamingFCLayer_Batch_5_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFCLayer_Batch_5_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFCLayer_Batch_5_out_V_V_TVALID),
        .weights_V_V_TDATA(StreamingFCLayer_Batch_5_wstrm_m_axis_0_TDATA),
        .weights_V_V_TREADY(StreamingFCLayer_Batch_5_wstrm_m_axis_0_TREADY),
        .weights_V_V_TVALID(StreamingFCLayer_Batch_5_wstrm_m_axis_0_TVALID));
  finn_design_StreamingFCLayer_Batch_5_wstrm_0 StreamingFCLayer_Batch_5_wstrm
       (.aclk(ap_clk_1),
        .araddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .aresetn(ap_rst_n_1),
        .arprot({1'b0,1'b0,1'b0}),
        .arvalid(1'b0),
        .awaddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .awprot({1'b0,1'b0,1'b0}),
        .awvalid(1'b0),
        .bready(1'b0),
        .m_axis_0_tdata(StreamingFCLayer_Batch_5_wstrm_m_axis_0_TDATA),
        .m_axis_0_tready(StreamingFCLayer_Batch_5_wstrm_m_axis_0_TREADY),
        .m_axis_0_tvalid(StreamingFCLayer_Batch_5_wstrm_m_axis_0_TVALID),
        .rready(1'b0),
        .wdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .wstrb({1'b1,1'b1,1'b1,1'b1}),
        .wvalid(1'b0));
endmodule

module StreamingFCLayer_Batch_6_imp_1Y3EON0
   (ap_clk,
    ap_rst_n,
    in0_V_V_tdata,
    in0_V_V_tready,
    in0_V_V_tvalid,
    out_V_V_tdata,
    out_V_V_tready,
    out_V_V_tvalid);
  input ap_clk;
  input ap_rst_n;
  input [7:0]in0_V_V_tdata;
  output in0_V_V_tready;
  input in0_V_V_tvalid;
  output [15:0]out_V_V_tdata;
  input out_V_V_tready;
  output out_V_V_tvalid;

  wire [15:0]StreamingFCLayer_Batch_6_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_6_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_6_out_V_V_TVALID;
  wire [7:0]StreamingFCLayer_Batch_6_wstrm_m_axis_0_TDATA;
  wire StreamingFCLayer_Batch_6_wstrm_m_axis_0_TREADY;
  wire StreamingFCLayer_Batch_6_wstrm_m_axis_0_TVALID;
  wire ap_clk_1;
  wire ap_rst_n_1;
  wire [7:0]in0_V_V_1_TDATA;
  wire in0_V_V_1_TREADY;
  wire in0_V_V_1_TVALID;

  assign StreamingFCLayer_Batch_6_out_V_V_TREADY = out_V_V_tready;
  assign ap_clk_1 = ap_clk;
  assign ap_rst_n_1 = ap_rst_n;
  assign in0_V_V_1_TDATA = in0_V_V_tdata[7:0];
  assign in0_V_V_1_TVALID = in0_V_V_tvalid;
  assign in0_V_V_tready = in0_V_V_1_TREADY;
  assign out_V_V_tdata[15:0] = StreamingFCLayer_Batch_6_out_V_V_TDATA;
  assign out_V_V_tvalid = StreamingFCLayer_Batch_6_out_V_V_TVALID;
  finn_design_StreamingFCLayer_Batch_6_0 StreamingFCLayer_Batch_6
       (.ap_clk(ap_clk_1),
        .ap_rst_n(ap_rst_n_1),
        .in0_V_V_TDATA(in0_V_V_1_TDATA),
        .in0_V_V_TREADY(in0_V_V_1_TREADY),
        .in0_V_V_TVALID(in0_V_V_1_TVALID),
        .out_V_V_TDATA(StreamingFCLayer_Batch_6_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFCLayer_Batch_6_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFCLayer_Batch_6_out_V_V_TVALID),
        .weights_V_V_TDATA(StreamingFCLayer_Batch_6_wstrm_m_axis_0_TDATA),
        .weights_V_V_TREADY(StreamingFCLayer_Batch_6_wstrm_m_axis_0_TREADY),
        .weights_V_V_TVALID(StreamingFCLayer_Batch_6_wstrm_m_axis_0_TVALID));
  finn_design_StreamingFCLayer_Batch_6_wstrm_0 StreamingFCLayer_Batch_6_wstrm
       (.aclk(ap_clk_1),
        .araddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .aresetn(ap_rst_n_1),
        .arprot({1'b0,1'b0,1'b0}),
        .arvalid(1'b0),
        .awaddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .awprot({1'b0,1'b0,1'b0}),
        .awvalid(1'b0),
        .bready(1'b0),
        .m_axis_0_tdata(StreamingFCLayer_Batch_6_wstrm_m_axis_0_TDATA),
        .m_axis_0_tready(StreamingFCLayer_Batch_6_wstrm_m_axis_0_TREADY),
        .m_axis_0_tvalid(StreamingFCLayer_Batch_6_wstrm_m_axis_0_TVALID),
        .rready(1'b0),
        .wdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .wstrb({1'b1,1'b1,1'b1,1'b1}),
        .wvalid(1'b0));
endmodule

(* CORE_GENERATION_INFO = "finn_design,IP_Integrator,{x_ipVendor=xilinx.com,x_ipLibrary=BlockDiagram,x_ipName=finn_design,x_ipVersion=1.00.a,x_ipLanguage=VERILOG,numBlks=55,numReposBlks=48,numNonXlnxBlks=0,numHierBlks=7,maxHierDepth=1,numSysgenBlks=0,numHlsBlks=21,numHdlrefBlks=0,numPkgbdBlks=0,bdsource=USER,synth_mode=OOC_per_IP}" *) (* HW_HANDOFF = "finn_design.hwdef" *) 
module finn_design
   (ap_clk,
    ap_rst_n,
    m_axis_0_tdata,
    m_axis_0_tready,
    m_axis_0_tvalid,
    m_axis_1_tdata,
    m_axis_1_tready,
    m_axis_1_tvalid,
    m_axis_2_tdata,
    m_axis_2_tready,
    m_axis_2_tvalid,
    s_axis_0_tdata,
    s_axis_0_tready,
    s_axis_0_tvalid,
    s_axis_1_tdata,
    s_axis_1_tready,
    s_axis_1_tvalid,
    s_axis_2_tdata,
    s_axis_2_tready,
    s_axis_2_tvalid);
  (* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 CLK.AP_CLK CLK" *) (* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME CLK.AP_CLK, ASSOCIATED_BUSIF s_axis_0:s_axis_1:s_axis_2:m_axis_0:m_axis_1:m_axis_2, ASSOCIATED_RESET ap_rst_n, CLK_DOMAIN finn_design_ap_clk_0, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, INSERT_VIP 0, PHASE 0.000" *) input ap_clk;
  (* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 RST.AP_RST_N RST" *) (* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME RST.AP_RST_N, INSERT_VIP 0, POLARITY ACTIVE_LOW" *) input ap_rst_n;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 " *) (* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME m_axis_0, CLK_DOMAIN finn_design_ap_clk_0, FREQ_HZ 100000000.000000, HAS_TKEEP 0, HAS_TLAST 0, HAS_TREADY 1, HAS_TSTRB 0, INSERT_VIP 0, LAYERED_METADATA undef, PHASE 0.000, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0" *) output [7:0]m_axis_0_tdata;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 " *) input m_axis_0_tready;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_0 " *) output m_axis_0_tvalid;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_1 " *) (* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME m_axis_1, CLK_DOMAIN finn_design_ap_clk_0, FREQ_HZ 100000000.000000, HAS_TKEEP 0, HAS_TLAST 0, HAS_TREADY 1, HAS_TSTRB 0, INSERT_VIP 0, LAYERED_METADATA undef, PHASE 0.000, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0" *) output [7:0]m_axis_1_tdata;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_1 " *) input m_axis_1_tready;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_1 " *) output m_axis_1_tvalid;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_2 " *) (* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME m_axis_2, CLK_DOMAIN finn_design_ap_clk_0, FREQ_HZ 100000000.000000, HAS_TKEEP 0, HAS_TLAST 0, HAS_TREADY 1, HAS_TSTRB 0, INSERT_VIP 0, LAYERED_METADATA undef, PHASE 0.000, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0" *) output [7:0]m_axis_2_tdata;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_2 " *) input m_axis_2_tready;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 m_axis_2 " *) output m_axis_2_tvalid;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 s_axis_0 " *) (* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axis_0, CLK_DOMAIN finn_design_ap_clk_0, FREQ_HZ 100000000.000000, HAS_TKEEP 0, HAS_TLAST 0, HAS_TREADY 1, HAS_TSTRB 0, INSERT_VIP 0, LAYERED_METADATA undef, PHASE 0.000, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0" *) input [7:0]s_axis_0_tdata;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 s_axis_0 " *) output s_axis_0_tready;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 s_axis_0 " *) input s_axis_0_tvalid;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 s_axis_1 " *) (* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axis_1, CLK_DOMAIN finn_design_ap_clk_0, FREQ_HZ 100000000.000000, HAS_TKEEP 0, HAS_TLAST 0, HAS_TREADY 1, HAS_TSTRB 0, INSERT_VIP 0, LAYERED_METADATA undef, PHASE 0.000, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0" *) input [7:0]s_axis_1_tdata;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 s_axis_1 " *) output s_axis_1_tready;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 s_axis_1 " *) input s_axis_1_tvalid;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 s_axis_2 " *) (* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axis_2, CLK_DOMAIN finn_design_ap_clk_0, FREQ_HZ 100000000.000000, HAS_TKEEP 0, HAS_TLAST 0, HAS_TREADY 1, HAS_TSTRB 0, INSERT_VIP 0, LAYERED_METADATA undef, PHASE 0.000, TDATA_NUM_BYTES 2, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0" *) input [15:0]s_axis_2_tdata;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 s_axis_2 " *) output s_axis_2_tready;
  (* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 s_axis_2 " *) input s_axis_2_tvalid;

  wire [7:0]ConvolutionInputGenerator_0_out_V_V_TDATA;
  wire ConvolutionInputGenerator_0_out_V_V_TREADY;
  wire ConvolutionInputGenerator_0_out_V_V_TVALID;
  wire [15:0]ConvolutionInputGenerator_1_out_V_V_TDATA;
  wire ConvolutionInputGenerator_1_out_V_V_TREADY;
  wire ConvolutionInputGenerator_1_out_V_V_TVALID;
  wire [23:0]ConvolutionInputGenerator_2_out_V_V_TDATA;
  wire ConvolutionInputGenerator_2_out_V_V_TREADY;
  wire ConvolutionInputGenerator_2_out_V_V_TVALID;
  wire [31:0]ConvolutionInputGenerator_3_out_V_V_TDATA;
  wire ConvolutionInputGenerator_3_out_V_V_TREADY;
  wire ConvolutionInputGenerator_3_out_V_V_TVALID;
  wire [7:0]LabelSelect_Batch_0_out_V_V_TDATA;
  wire LabelSelect_Batch_0_out_V_V_TREADY;
  wire LabelSelect_Batch_0_out_V_V_TVALID;
  wire [23:0]StreamingDataWidthConverter_Batch_0_out_V_V_TDATA;
  wire StreamingDataWidthConverter_Batch_0_out_V_V_TREADY;
  wire StreamingDataWidthConverter_Batch_0_out_V_V_TVALID;
  wire [23:0]StreamingDataWidthConverter_Batch_1_out_V_V_TDATA;
  wire StreamingDataWidthConverter_Batch_1_out_V_V_TREADY;
  wire StreamingDataWidthConverter_Batch_1_out_V_V_TVALID;
  wire [31:0]StreamingDataWidthConverter_Batch_2_out_V_V_TDATA;
  wire StreamingDataWidthConverter_Batch_2_out_V_V_TREADY;
  wire StreamingDataWidthConverter_Batch_2_out_V_V_TVALID;
  wire [31:0]StreamingDataWidthConverter_Batch_3_out_V_V_TDATA;
  wire StreamingDataWidthConverter_Batch_3_out_V_V_TREADY;
  wire StreamingDataWidthConverter_Batch_3_out_V_V_TVALID;
  wire [31:0]StreamingDataWidthConverter_Batch_4_out_V_V_TDATA;
  wire StreamingDataWidthConverter_Batch_4_out_V_V_TREADY;
  wire StreamingDataWidthConverter_Batch_4_out_V_V_TVALID;
  wire [7:0]StreamingDataWidthConverter_Batch_5_out_V_V_TDATA;
  wire StreamingDataWidthConverter_Batch_5_out_V_V_TREADY;
  wire StreamingDataWidthConverter_Batch_5_out_V_V_TVALID;
  wire [95:0]StreamingFCLayer_Batch_0_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_0_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_0_out_V_V_TVALID;
  wire [15:0]StreamingFCLayer_Batch_1_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_1_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_1_out_V_V_TVALID;
  wire [15:0]StreamingFCLayer_Batch_2_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_2_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_2_out_V_V_TVALID;
  wire [15:0]StreamingFCLayer_Batch_3_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_3_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_3_out_V_V_TVALID;
  wire [15:0]StreamingFCLayer_Batch_4_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_4_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_4_out_V_V_TVALID;
  wire [15:0]StreamingFCLayer_Batch_5_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_5_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_5_out_V_V_TVALID;
  wire [15:0]StreamingFCLayer_Batch_6_out_V_V_TDATA;
  wire StreamingFCLayer_Batch_6_out_V_V_TREADY;
  wire StreamingFCLayer_Batch_6_out_V_V_TVALID;
  wire [7:0]StreamingFIFO_0_out_V_V_TDATA;
  wire StreamingFIFO_0_out_V_V_TREADY;
  wire StreamingFIFO_0_out_V_V_TVALID;
  wire [15:0]StreamingFIFO_10_out_V_V_TDATA;
  wire StreamingFIFO_10_out_V_V_TREADY;
  wire StreamingFIFO_10_out_V_V_TVALID;
  wire [15:0]StreamingFIFO_11_out_V_V_TDATA;
  wire StreamingFIFO_11_out_V_V_TREADY;
  wire StreamingFIFO_11_out_V_V_TVALID;
  wire [31:0]StreamingFIFO_12_out_V_V_TDATA;
  wire StreamingFIFO_12_out_V_V_TREADY;
  wire StreamingFIFO_12_out_V_V_TVALID;
  wire [31:0]StreamingFIFO_13_out_V_V_TDATA;
  wire StreamingFIFO_13_out_V_V_TREADY;
  wire StreamingFIFO_13_out_V_V_TVALID;
  wire [15:0]StreamingFIFO_14_out_V_V_TDATA;
  wire StreamingFIFO_14_out_V_V_TREADY;
  wire StreamingFIFO_14_out_V_V_TVALID;
  wire [31:0]StreamingFIFO_15_out_V_V_TDATA;
  wire StreamingFIFO_15_out_V_V_TREADY;
  wire StreamingFIFO_15_out_V_V_TVALID;
  wire [7:0]StreamingFIFO_16_out_V_V_TDATA;
  wire StreamingFIFO_16_out_V_V_TREADY;
  wire StreamingFIFO_16_out_V_V_TVALID;
  wire [15:0]StreamingFIFO_17_out_V_V_TDATA;
  wire StreamingFIFO_17_out_V_V_TREADY;
  wire StreamingFIFO_17_out_V_V_TVALID;
  wire [15:0]StreamingFIFO_18_out_V_V_TDATA;
  wire StreamingFIFO_18_out_V_V_TREADY;
  wire StreamingFIFO_18_out_V_V_TVALID;
  wire [7:0]StreamingFIFO_19_out_V_V_TDATA;
  wire StreamingFIFO_19_out_V_V_TREADY;
  wire StreamingFIFO_19_out_V_V_TVALID;
  wire [7:0]StreamingFIFO_1_out_V_V_TDATA;
  wire StreamingFIFO_1_out_V_V_TREADY;
  wire StreamingFIFO_1_out_V_V_TVALID;
  wire [15:0]StreamingFIFO_2_out_V_V_TDATA;
  wire StreamingFIFO_2_out_V_V_TREADY;
  wire StreamingFIFO_2_out_V_V_TVALID;
  wire [7:0]StreamingFIFO_3_out_V_V_TDATA;
  wire StreamingFIFO_3_out_V_V_TREADY;
  wire StreamingFIFO_3_out_V_V_TVALID;
  wire [95:0]StreamingFIFO_4_out_V_V_TDATA;
  wire StreamingFIFO_4_out_V_V_TREADY;
  wire StreamingFIFO_4_out_V_V_TVALID;
  wire [15:0]StreamingFIFO_5_out_V_V_TDATA;
  wire StreamingFIFO_5_out_V_V_TREADY;
  wire StreamingFIFO_5_out_V_V_TVALID;
  wire [23:0]StreamingFIFO_6_out_V_V_TDATA;
  wire StreamingFIFO_6_out_V_V_TREADY;
  wire StreamingFIFO_6_out_V_V_TVALID;
  wire [23:0]StreamingFIFO_7_out_V_V_TDATA;
  wire StreamingFIFO_7_out_V_V_TREADY;
  wire StreamingFIFO_7_out_V_V_TVALID;
  wire [31:0]StreamingFIFO_8_out_V_V_TDATA;
  wire StreamingFIFO_8_out_V_V_TREADY;
  wire StreamingFIFO_8_out_V_V_TVALID;
  wire [23:0]StreamingFIFO_9_out_V_V_TDATA;
  wire StreamingFIFO_9_out_V_V_TREADY;
  wire StreamingFIFO_9_out_V_V_TVALID;
  wire [7:0]Thresholding_Batch_0_out_V_V_TDATA;
  wire Thresholding_Batch_0_out_V_V_TREADY;
  wire Thresholding_Batch_0_out_V_V_TVALID;
  wire [7:0]Thresholding_Batch_1_out_V_V_TDATA;
  wire Thresholding_Batch_1_out_V_V_TREADY;
  wire Thresholding_Batch_1_out_V_V_TVALID;
  wire [7:0]Thresholding_Batch_2_out_V_V_TDATA;
  wire Thresholding_Batch_2_out_V_V_TREADY;
  wire Thresholding_Batch_2_out_V_V_TVALID;
  wire ap_clk_0_1;
  wire ap_rst_n_0_1;
  wire [7:0]in0_V_V_0_1_TDATA;
  wire in0_V_V_0_1_TREADY;
  wire in0_V_V_0_1_TVALID;
  wire [7:0]in0_V_V_0_2_TDATA;
  wire in0_V_V_0_2_TREADY;
  wire in0_V_V_0_2_TVALID;
  wire [15:0]in0_V_V_0_3_TDATA;
  wire in0_V_V_0_3_TREADY;
  wire in0_V_V_0_3_TVALID;

  assign StreamingFIFO_19_out_V_V_TREADY = m_axis_2_tready;
  assign Thresholding_Batch_1_out_V_V_TREADY = m_axis_0_tready;
  assign Thresholding_Batch_2_out_V_V_TREADY = m_axis_1_tready;
  assign ap_clk_0_1 = ap_clk;
  assign ap_rst_n_0_1 = ap_rst_n;
  assign in0_V_V_0_1_TDATA = s_axis_0_tdata[7:0];
  assign in0_V_V_0_1_TVALID = s_axis_0_tvalid;
  assign in0_V_V_0_2_TDATA = s_axis_1_tdata[7:0];
  assign in0_V_V_0_2_TVALID = s_axis_1_tvalid;
  assign in0_V_V_0_3_TDATA = s_axis_2_tdata[15:0];
  assign in0_V_V_0_3_TVALID = s_axis_2_tvalid;
  assign m_axis_0_tdata[7:0] = Thresholding_Batch_1_out_V_V_TDATA;
  assign m_axis_0_tvalid = Thresholding_Batch_1_out_V_V_TVALID;
  assign m_axis_1_tdata[7:0] = Thresholding_Batch_2_out_V_V_TDATA;
  assign m_axis_1_tvalid = Thresholding_Batch_2_out_V_V_TVALID;
  assign m_axis_2_tdata[7:0] = StreamingFIFO_19_out_V_V_TDATA;
  assign m_axis_2_tvalid = StreamingFIFO_19_out_V_V_TVALID;
  assign s_axis_0_tready = in0_V_V_0_1_TREADY;
  assign s_axis_1_tready = in0_V_V_0_2_TREADY;
  assign s_axis_2_tready = in0_V_V_0_3_TREADY;
  finn_design_ConvolutionInputGenerator_0_0 ConvolutionInputGenerator_0
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(in0_V_V_0_2_TDATA),
        .in0_V_V_TREADY(in0_V_V_0_2_TREADY),
        .in0_V_V_TVALID(in0_V_V_0_2_TVALID),
        .out_V_V_TDATA(ConvolutionInputGenerator_0_out_V_V_TDATA),
        .out_V_V_TREADY(ConvolutionInputGenerator_0_out_V_V_TREADY),
        .out_V_V_TVALID(ConvolutionInputGenerator_0_out_V_V_TVALID));
  finn_design_ConvolutionInputGenerator_1_0 ConvolutionInputGenerator_1
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(in0_V_V_0_3_TDATA),
        .in0_V_V_TREADY(in0_V_V_0_3_TREADY),
        .in0_V_V_TVALID(in0_V_V_0_3_TVALID),
        .out_V_V_TDATA(ConvolutionInputGenerator_1_out_V_V_TDATA),
        .out_V_V_TREADY(ConvolutionInputGenerator_1_out_V_V_TREADY),
        .out_V_V_TVALID(ConvolutionInputGenerator_1_out_V_V_TVALID));
  finn_design_ConvolutionInputGenerator_2_0 ConvolutionInputGenerator_2
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_6_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_6_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_6_out_V_V_TVALID),
        .out_V_V_TDATA(ConvolutionInputGenerator_2_out_V_V_TDATA),
        .out_V_V_TREADY(ConvolutionInputGenerator_2_out_V_V_TREADY),
        .out_V_V_TVALID(ConvolutionInputGenerator_2_out_V_V_TVALID));
  finn_design_ConvolutionInputGenerator_3_0 ConvolutionInputGenerator_3
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_13_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_13_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_13_out_V_V_TVALID),
        .out_V_V_TDATA(ConvolutionInputGenerator_3_out_V_V_TDATA),
        .out_V_V_TREADY(ConvolutionInputGenerator_3_out_V_V_TREADY),
        .out_V_V_TVALID(ConvolutionInputGenerator_3_out_V_V_TVALID));
  finn_design_LabelSelect_Batch_0_0 LabelSelect_Batch_0
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_18_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_18_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_18_out_V_V_TVALID),
        .out_V_V_TDATA(LabelSelect_Batch_0_out_V_V_TDATA),
        .out_V_V_TREADY(LabelSelect_Batch_0_out_V_V_TREADY),
        .out_V_V_TVALID(LabelSelect_Batch_0_out_V_V_TVALID));
  finn_design_StreamingDataWidthConverter_Batch_0_0 StreamingDataWidthConverter_Batch_0
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_3_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_3_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_3_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingDataWidthConverter_Batch_0_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingDataWidthConverter_Batch_0_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingDataWidthConverter_Batch_0_out_V_V_TVALID));
  finn_design_StreamingDataWidthConverter_Batch_1_0 StreamingDataWidthConverter_Batch_1
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_4_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_4_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_4_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingDataWidthConverter_Batch_1_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingDataWidthConverter_Batch_1_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingDataWidthConverter_Batch_1_out_V_V_TVALID));
  finn_design_StreamingDataWidthConverter_Batch_2_0 StreamingDataWidthConverter_Batch_2
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_5_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_5_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_5_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingDataWidthConverter_Batch_2_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingDataWidthConverter_Batch_2_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingDataWidthConverter_Batch_2_out_V_V_TVALID));
  finn_design_StreamingDataWidthConverter_Batch_3_0 StreamingDataWidthConverter_Batch_3
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_10_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_10_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_10_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingDataWidthConverter_Batch_3_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingDataWidthConverter_Batch_3_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingDataWidthConverter_Batch_3_out_V_V_TVALID));
  finn_design_StreamingDataWidthConverter_Batch_4_0 StreamingDataWidthConverter_Batch_4
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_11_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_11_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_11_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingDataWidthConverter_Batch_4_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingDataWidthConverter_Batch_4_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingDataWidthConverter_Batch_4_out_V_V_TVALID));
  finn_design_StreamingDataWidthConverter_Batch_5_0 StreamingDataWidthConverter_Batch_5
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_14_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_14_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_14_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingDataWidthConverter_Batch_5_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingDataWidthConverter_Batch_5_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingDataWidthConverter_Batch_5_out_V_V_TVALID));
  StreamingFCLayer_Batch_0_imp_5FXKV0 StreamingFCLayer_Batch_0
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_tdata(StreamingFIFO_1_out_V_V_TDATA),
        .in0_V_V_tready(StreamingFIFO_1_out_V_V_TREADY),
        .in0_V_V_tvalid(StreamingFIFO_1_out_V_V_TVALID),
        .out_V_V_tdata(StreamingFCLayer_Batch_0_out_V_V_TDATA),
        .out_V_V_tready(StreamingFCLayer_Batch_0_out_V_V_TREADY),
        .out_V_V_tvalid(StreamingFCLayer_Batch_0_out_V_V_TVALID));
  StreamingFCLayer_Batch_1_imp_11SOJ3N StreamingFCLayer_Batch_1
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_tdata(StreamingFIFO_2_out_V_V_TDATA),
        .in0_V_V_tready(StreamingFIFO_2_out_V_V_TREADY),
        .in0_V_V_tvalid(StreamingFIFO_2_out_V_V_TVALID),
        .out_V_V_tdata(StreamingFCLayer_Batch_1_out_V_V_TDATA),
        .out_V_V_tready(StreamingFCLayer_Batch_1_out_V_V_TREADY),
        .out_V_V_tvalid(StreamingFCLayer_Batch_1_out_V_V_TVALID));
  StreamingFCLayer_Batch_2_imp_1YXLQV7 StreamingFCLayer_Batch_2
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_tdata(StreamingFIFO_8_out_V_V_TDATA),
        .in0_V_V_tready(StreamingFIFO_8_out_V_V_TREADY),
        .in0_V_V_tvalid(StreamingFIFO_8_out_V_V_TVALID),
        .out_V_V_tdata(StreamingFCLayer_Batch_2_out_V_V_TDATA),
        .out_V_V_tready(StreamingFCLayer_Batch_2_out_V_V_TREADY),
        .out_V_V_tvalid(StreamingFCLayer_Batch_2_out_V_V_TVALID));
  StreamingFCLayer_Batch_3_imp_RR03E4 StreamingFCLayer_Batch_3
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_tdata(StreamingFIFO_9_out_V_V_TDATA),
        .in0_V_V_tready(StreamingFIFO_9_out_V_V_TREADY),
        .in0_V_V_tvalid(StreamingFIFO_9_out_V_V_TVALID),
        .out_V_V_tdata(StreamingFCLayer_Batch_3_out_V_V_TDATA),
        .out_V_V_tready(StreamingFCLayer_Batch_3_out_V_V_TREADY),
        .out_V_V_tvalid(StreamingFCLayer_Batch_3_out_V_V_TVALID));
  StreamingFCLayer_Batch_4_imp_4LW78J StreamingFCLayer_Batch_4
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_tdata(StreamingFIFO_12_out_V_V_TDATA),
        .in0_V_V_tready(StreamingFIFO_12_out_V_V_TREADY),
        .in0_V_V_tvalid(StreamingFIFO_12_out_V_V_TVALID),
        .out_V_V_tdata(StreamingFCLayer_Batch_4_out_V_V_TDATA),
        .out_V_V_tready(StreamingFCLayer_Batch_4_out_V_V_TREADY),
        .out_V_V_tvalid(StreamingFCLayer_Batch_4_out_V_V_TVALID));
  StreamingFCLayer_Batch_5_imp_12MW1JG StreamingFCLayer_Batch_5
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_tdata(StreamingFIFO_15_out_V_V_TDATA),
        .in0_V_V_tready(StreamingFIFO_15_out_V_V_TREADY),
        .in0_V_V_tvalid(StreamingFIFO_15_out_V_V_TVALID),
        .out_V_V_tdata(StreamingFCLayer_Batch_5_out_V_V_TDATA),
        .out_V_V_tready(StreamingFCLayer_Batch_5_out_V_V_TREADY),
        .out_V_V_tvalid(StreamingFCLayer_Batch_5_out_V_V_TVALID));
  StreamingFCLayer_Batch_6_imp_1Y3EON0 StreamingFCLayer_Batch_6
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_tdata(StreamingFIFO_16_out_V_V_TDATA),
        .in0_V_V_tready(StreamingFIFO_16_out_V_V_TREADY),
        .in0_V_V_tvalid(StreamingFIFO_16_out_V_V_TVALID),
        .out_V_V_tdata(StreamingFCLayer_Batch_6_out_V_V_TDATA),
        .out_V_V_tready(StreamingFCLayer_Batch_6_out_V_V_TREADY),
        .out_V_V_tvalid(StreamingFCLayer_Batch_6_out_V_V_TVALID));
  finn_design_StreamingFIFO_0_0 StreamingFIFO_0
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(in0_V_V_0_1_TDATA),
        .in0_V_V_TREADY(in0_V_V_0_1_TREADY),
        .in0_V_V_TVALID(in0_V_V_0_1_TVALID),
        .out_V_V_TDATA(StreamingFIFO_0_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_0_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_0_out_V_V_TVALID));
  finn_design_StreamingFIFO_1_0 StreamingFIFO_1
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(ConvolutionInputGenerator_0_out_V_V_TDATA),
        .in0_V_V_TREADY(ConvolutionInputGenerator_0_out_V_V_TREADY),
        .in0_V_V_TVALID(ConvolutionInputGenerator_0_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_1_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_1_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_1_out_V_V_TVALID));
  finn_design_StreamingFIFO_10_0 StreamingFIFO_10
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFCLayer_Batch_2_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFCLayer_Batch_2_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFCLayer_Batch_2_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_10_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_10_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_10_out_V_V_TVALID));
  finn_design_StreamingFIFO_11_0 StreamingFIFO_11
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFCLayer_Batch_3_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFCLayer_Batch_3_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFCLayer_Batch_3_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_11_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_11_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_11_out_V_V_TVALID));
  finn_design_StreamingFIFO_12_0 StreamingFIFO_12
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingDataWidthConverter_Batch_3_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingDataWidthConverter_Batch_3_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingDataWidthConverter_Batch_3_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_12_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_12_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_12_out_V_V_TVALID));
  finn_design_StreamingFIFO_13_0 StreamingFIFO_13
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingDataWidthConverter_Batch_4_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingDataWidthConverter_Batch_4_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingDataWidthConverter_Batch_4_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_13_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_13_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_13_out_V_V_TVALID));
  finn_design_StreamingFIFO_14_0 StreamingFIFO_14
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFCLayer_Batch_4_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFCLayer_Batch_4_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFCLayer_Batch_4_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_14_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_14_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_14_out_V_V_TVALID));
  finn_design_StreamingFIFO_15_0 StreamingFIFO_15
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(ConvolutionInputGenerator_3_out_V_V_TDATA),
        .in0_V_V_TREADY(ConvolutionInputGenerator_3_out_V_V_TREADY),
        .in0_V_V_TVALID(ConvolutionInputGenerator_3_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_15_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_15_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_15_out_V_V_TVALID));
  finn_design_StreamingFIFO_16_0 StreamingFIFO_16
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingDataWidthConverter_Batch_5_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingDataWidthConverter_Batch_5_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingDataWidthConverter_Batch_5_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_16_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_16_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_16_out_V_V_TVALID));
  finn_design_StreamingFIFO_17_0 StreamingFIFO_17
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFCLayer_Batch_5_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFCLayer_Batch_5_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFCLayer_Batch_5_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_17_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_17_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_17_out_V_V_TVALID));
  finn_design_StreamingFIFO_18_0 StreamingFIFO_18
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFCLayer_Batch_6_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFCLayer_Batch_6_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFCLayer_Batch_6_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_18_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_18_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_18_out_V_V_TVALID));
  finn_design_StreamingFIFO_19_0 StreamingFIFO_19
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(LabelSelect_Batch_0_out_V_V_TDATA),
        .in0_V_V_TREADY(LabelSelect_Batch_0_out_V_V_TREADY),
        .in0_V_V_TVALID(LabelSelect_Batch_0_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_19_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_19_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_19_out_V_V_TVALID));
  finn_design_StreamingFIFO_2_0 StreamingFIFO_2
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(ConvolutionInputGenerator_1_out_V_V_TDATA),
        .in0_V_V_TREADY(ConvolutionInputGenerator_1_out_V_V_TREADY),
        .in0_V_V_TVALID(ConvolutionInputGenerator_1_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_2_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_2_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_2_out_V_V_TVALID));
  finn_design_StreamingFIFO_3_0 StreamingFIFO_3
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(Thresholding_Batch_0_out_V_V_TDATA),
        .in0_V_V_TREADY(Thresholding_Batch_0_out_V_V_TREADY),
        .in0_V_V_TVALID(Thresholding_Batch_0_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_3_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_3_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_3_out_V_V_TVALID));
  finn_design_StreamingFIFO_4_0 StreamingFIFO_4
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFCLayer_Batch_0_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFCLayer_Batch_0_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFCLayer_Batch_0_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_4_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_4_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_4_out_V_V_TVALID));
  finn_design_StreamingFIFO_5_0 StreamingFIFO_5
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFCLayer_Batch_1_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFCLayer_Batch_1_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFCLayer_Batch_1_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_5_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_5_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_5_out_V_V_TVALID));
  finn_design_StreamingFIFO_6_0 StreamingFIFO_6
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingDataWidthConverter_Batch_0_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingDataWidthConverter_Batch_0_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingDataWidthConverter_Batch_0_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_6_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_6_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_6_out_V_V_TVALID));
  finn_design_StreamingFIFO_7_0 StreamingFIFO_7
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingDataWidthConverter_Batch_1_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingDataWidthConverter_Batch_1_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingDataWidthConverter_Batch_1_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_7_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_7_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_7_out_V_V_TVALID));
  finn_design_StreamingFIFO_8_0 StreamingFIFO_8
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingDataWidthConverter_Batch_2_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingDataWidthConverter_Batch_2_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingDataWidthConverter_Batch_2_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_8_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_8_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_8_out_V_V_TVALID));
  finn_design_StreamingFIFO_9_0 StreamingFIFO_9
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(ConvolutionInputGenerator_2_out_V_V_TDATA),
        .in0_V_V_TREADY(ConvolutionInputGenerator_2_out_V_V_TREADY),
        .in0_V_V_TVALID(ConvolutionInputGenerator_2_out_V_V_TVALID),
        .out_V_V_TDATA(StreamingFIFO_9_out_V_V_TDATA),
        .out_V_V_TREADY(StreamingFIFO_9_out_V_V_TREADY),
        .out_V_V_TVALID(StreamingFIFO_9_out_V_V_TVALID));
  finn_design_Thresholding_Batch_0_0 Thresholding_Batch_0
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_0_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_0_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_0_out_V_V_TVALID),
        .out_V_V_TDATA(Thresholding_Batch_0_out_V_V_TDATA),
        .out_V_V_TREADY(Thresholding_Batch_0_out_V_V_TREADY),
        .out_V_V_TVALID(Thresholding_Batch_0_out_V_V_TVALID));
  finn_design_Thresholding_Batch_1_0 Thresholding_Batch_1
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_7_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_7_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_7_out_V_V_TVALID),
        .out_V_V_TDATA(Thresholding_Batch_1_out_V_V_TDATA),
        .out_V_V_TREADY(Thresholding_Batch_1_out_V_V_TREADY),
        .out_V_V_TVALID(Thresholding_Batch_1_out_V_V_TVALID));
  finn_design_Thresholding_Batch_2_0 Thresholding_Batch_2
       (.ap_clk(ap_clk_0_1),
        .ap_rst_n(ap_rst_n_0_1),
        .in0_V_V_TDATA(StreamingFIFO_17_out_V_V_TDATA),
        .in0_V_V_TREADY(StreamingFIFO_17_out_V_V_TREADY),
        .in0_V_V_TVALID(StreamingFIFO_17_out_V_V_TVALID),
        .out_V_V_TDATA(Thresholding_Batch_2_out_V_V_TDATA),
        .out_V_V_TREADY(Thresholding_Batch_2_out_V_V_TREADY),
        .out_V_V_TVALID(Thresholding_Batch_2_out_V_V_TVALID));
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActPgM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActPgM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActPgM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActPgM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActPgM_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActPgM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/bc91/hdl/verilog/StreamingFCLayer_Batch_6_StreamingFCLayer_bkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module StreamingFCLayer_Batch_6_StreamingFCLayer_bkb #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH       = 32,
    din5_WIDTH       = 32,
    din6_WIDTH       = 32,
    din7_WIDTH       = 32,
    din8_WIDTH       = 32,
    din9_WIDTH       = 32,
    din10_WIDTH       = 32,
    din11_WIDTH       = 32,
    din12_WIDTH       = 32,
    din13_WIDTH       = 32,
    din14_WIDTH       = 32,
    din15_WIDTH       = 32,
    din16_WIDTH       = 32,
    din17_WIDTH       = 32,
    din18_WIDTH       = 32,
    din19_WIDTH       = 32,
    din20_WIDTH       = 32,
    din21_WIDTH       = 32,
    din22_WIDTH       = 32,
    din23_WIDTH       = 32,
    din24_WIDTH       = 32,
    din25_WIDTH       = 32,
    din26_WIDTH       = 32,
    din27_WIDTH       = 32,
    din28_WIDTH       = 32,
    din29_WIDTH       = 32,
    din30_WIDTH       = 32,
    din31_WIDTH       = 32,
    din32_WIDTH       = 32,
    din33_WIDTH       = 32,
    din34_WIDTH       = 32,
    din35_WIDTH       = 32,
    din36_WIDTH       = 32,
    din37_WIDTH       = 32,
    din38_WIDTH       = 32,
    din39_WIDTH       = 32,
    din40_WIDTH       = 32,
    din41_WIDTH       = 32,
    din42_WIDTH       = 32,
    din43_WIDTH       = 32,
    din44_WIDTH       = 32,
    din45_WIDTH       = 32,
    din46_WIDTH       = 32,
    din47_WIDTH       = 32,
    din48_WIDTH       = 32,
    din49_WIDTH       = 32,
    din50_WIDTH       = 32,
    din51_WIDTH       = 32,
    din52_WIDTH       = 32,
    din53_WIDTH       = 32,
    din54_WIDTH       = 32,
    din55_WIDTH       = 32,
    din56_WIDTH       = 32,
    din57_WIDTH       = 32,
    din58_WIDTH       = 32,
    din59_WIDTH       = 32,
    din60_WIDTH       = 32,
    din61_WIDTH       = 32,
    din62_WIDTH       = 32,
    din63_WIDTH       = 32,
    din64_WIDTH       = 32,
    din65_WIDTH       = 32,
    din66_WIDTH       = 32,
    din67_WIDTH       = 32,
    din68_WIDTH       = 32,
    din69_WIDTH       = 32,
    din70_WIDTH       = 32,
    din71_WIDTH       = 32,
    din72_WIDTH       = 32,
    din73_WIDTH       = 32,
    din74_WIDTH       = 32,
    din75_WIDTH       = 32,
    din76_WIDTH       = 32,
    din77_WIDTH       = 32,
    din78_WIDTH       = 32,
    din79_WIDTH       = 32,
    din80_WIDTH       = 32,
    din81_WIDTH       = 32,
    din82_WIDTH       = 32,
    din83_WIDTH       = 32,
    din84_WIDTH       = 32,
    din85_WIDTH       = 32,
    din86_WIDTH       = 32,
    din87_WIDTH       = 32,
    din88_WIDTH       = 32,
    din89_WIDTH       = 32,
    din90_WIDTH       = 32,
    din91_WIDTH       = 32,
    din92_WIDTH       = 32,
    din93_WIDTH       = 32,
    din94_WIDTH       = 32,
    din95_WIDTH       = 32,
    din96_WIDTH       = 32,
    din97_WIDTH       = 32,
    din98_WIDTH       = 32,
    din99_WIDTH       = 32,
    din100_WIDTH       = 32,
    din101_WIDTH       = 32,
    din102_WIDTH       = 32,
    din103_WIDTH       = 32,
    din104_WIDTH       = 32,
    din105_WIDTH       = 32,
    din106_WIDTH       = 32,
    din107_WIDTH       = 32,
    din108_WIDTH       = 32,
    din109_WIDTH       = 32,
    din110_WIDTH       = 32,
    din111_WIDTH       = 32,
    din112_WIDTH       = 32,
    din113_WIDTH       = 32,
    din114_WIDTH       = 32,
    din115_WIDTH       = 32,
    din116_WIDTH       = 32,
    din117_WIDTH       = 32,
    din118_WIDTH       = 32,
    din119_WIDTH       = 32,
    din120_WIDTH       = 32,
    din121_WIDTH       = 32,
    din122_WIDTH       = 32,
    din123_WIDTH       = 32,
    din124_WIDTH       = 32,
    din125_WIDTH       = 32,
    din126_WIDTH       = 32,
    din127_WIDTH       = 32,
    din128_WIDTH       = 32,
    din129_WIDTH       = 32,
    din130_WIDTH       = 32,
    din131_WIDTH       = 32,
    din132_WIDTH       = 32,
    din133_WIDTH       = 32,
    din134_WIDTH       = 32,
    din135_WIDTH       = 32,
    din136_WIDTH       = 32,
    din137_WIDTH       = 32,
    din138_WIDTH       = 32,
    din139_WIDTH       = 32,
    din140_WIDTH       = 32,
    din141_WIDTH       = 32,
    din142_WIDTH       = 32,
    din143_WIDTH       = 32,
    din144_WIDTH       = 32,
    din145_WIDTH       = 32,
    din146_WIDTH       = 32,
    din147_WIDTH       = 32,
    din148_WIDTH       = 32,
    din149_WIDTH       = 32,
    din150_WIDTH       = 32,
    din151_WIDTH       = 32,
    din152_WIDTH       = 32,
    din153_WIDTH       = 32,
    din154_WIDTH       = 32,
    din155_WIDTH       = 32,
    din156_WIDTH       = 32,
    din157_WIDTH       = 32,
    din158_WIDTH       = 32,
    din159_WIDTH       = 32,
    din160_WIDTH       = 32,
    din161_WIDTH       = 32,
    din162_WIDTH       = 32,
    din163_WIDTH       = 32,
    din164_WIDTH       = 32,
    din165_WIDTH       = 32,
    din166_WIDTH       = 32,
    din167_WIDTH       = 32,
    din168_WIDTH       = 32,
    din169_WIDTH       = 32,
    din170_WIDTH       = 32,
    din171_WIDTH       = 32,
    din172_WIDTH       = 32,
    din173_WIDTH       = 32,
    din174_WIDTH       = 32,
    din175_WIDTH       = 32,
    din176_WIDTH       = 32,
    din177_WIDTH       = 32,
    din178_WIDTH       = 32,
    din179_WIDTH       = 32,
    din180_WIDTH       = 32,
    din181_WIDTH       = 32,
    din182_WIDTH       = 32,
    din183_WIDTH       = 32,
    din184_WIDTH       = 32,
    din185_WIDTH       = 32,
    din186_WIDTH       = 32,
    din187_WIDTH       = 32,
    din188_WIDTH       = 32,
    din189_WIDTH       = 32,
    din190_WIDTH       = 32,
    din191_WIDTH       = 32,
    din192_WIDTH       = 32,
    din193_WIDTH       = 32,
    din194_WIDTH       = 32,
    din195_WIDTH       = 32,
    din196_WIDTH       = 32,
    din197_WIDTH       = 32,
    din198_WIDTH       = 32,
    din199_WIDTH       = 32,
    din200_WIDTH       = 32,
    din201_WIDTH       = 32,
    din202_WIDTH       = 32,
    din203_WIDTH       = 32,
    din204_WIDTH       = 32,
    din205_WIDTH       = 32,
    din206_WIDTH       = 32,
    din207_WIDTH       = 32,
    din208_WIDTH       = 32,
    din209_WIDTH       = 32,
    din210_WIDTH       = 32,
    din211_WIDTH       = 32,
    din212_WIDTH       = 32,
    din213_WIDTH       = 32,
    din214_WIDTH       = 32,
    din215_WIDTH       = 32,
    din216_WIDTH       = 32,
    din217_WIDTH       = 32,
    din218_WIDTH       = 32,
    din219_WIDTH       = 32,
    din220_WIDTH       = 32,
    din221_WIDTH       = 32,
    din222_WIDTH       = 32,
    din223_WIDTH       = 32,
    din224_WIDTH       = 32,
    din225_WIDTH       = 32,
    din226_WIDTH       = 32,
    din227_WIDTH       = 32,
    din228_WIDTH       = 32,
    din229_WIDTH       = 32,
    din230_WIDTH       = 32,
    din231_WIDTH       = 32,
    din232_WIDTH       = 32,
    din233_WIDTH       = 32,
    din234_WIDTH       = 32,
    din235_WIDTH       = 32,
    din236_WIDTH       = 32,
    din237_WIDTH       = 32,
    din238_WIDTH       = 32,
    din239_WIDTH       = 32,
    din240_WIDTH       = 32,
    din241_WIDTH       = 32,
    din242_WIDTH       = 32,
    din243_WIDTH       = 32,
    din244_WIDTH       = 32,
    din245_WIDTH       = 32,
    din246_WIDTH       = 32,
    din247_WIDTH       = 32,
    din248_WIDTH       = 32,
    din249_WIDTH       = 32,
    din250_WIDTH       = 32,
    din251_WIDTH       = 32,
    din252_WIDTH       = 32,
    din253_WIDTH       = 32,
    din254_WIDTH       = 32,
    din255_WIDTH       = 32,
    din256_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [7 : 0]     din0,
    input  [7 : 0]     din1,
    input  [7 : 0]     din2,
    input  [7 : 0]     din3,
    input  [7 : 0]     din4,
    input  [7 : 0]     din5,
    input  [7 : 0]     din6,
    input  [7 : 0]     din7,
    input  [7 : 0]     din8,
    input  [7 : 0]     din9,
    input  [7 : 0]     din10,
    input  [7 : 0]     din11,
    input  [7 : 0]     din12,
    input  [7 : 0]     din13,
    input  [7 : 0]     din14,
    input  [7 : 0]     din15,
    input  [7 : 0]     din16,
    input  [7 : 0]     din17,
    input  [7 : 0]     din18,
    input  [7 : 0]     din19,
    input  [7 : 0]     din20,
    input  [7 : 0]     din21,
    input  [7 : 0]     din22,
    input  [7 : 0]     din23,
    input  [7 : 0]     din24,
    input  [7 : 0]     din25,
    input  [7 : 0]     din26,
    input  [7 : 0]     din27,
    input  [7 : 0]     din28,
    input  [7 : 0]     din29,
    input  [7 : 0]     din30,
    input  [7 : 0]     din31,
    input  [7 : 0]     din32,
    input  [7 : 0]     din33,
    input  [7 : 0]     din34,
    input  [7 : 0]     din35,
    input  [7 : 0]     din36,
    input  [7 : 0]     din37,
    input  [7 : 0]     din38,
    input  [7 : 0]     din39,
    input  [7 : 0]     din40,
    input  [7 : 0]     din41,
    input  [7 : 0]     din42,
    input  [7 : 0]     din43,
    input  [7 : 0]     din44,
    input  [7 : 0]     din45,
    input  [7 : 0]     din46,
    input  [7 : 0]     din47,
    input  [7 : 0]     din48,
    input  [7 : 0]     din49,
    input  [7 : 0]     din50,
    input  [7 : 0]     din51,
    input  [7 : 0]     din52,
    input  [7 : 0]     din53,
    input  [7 : 0]     din54,
    input  [7 : 0]     din55,
    input  [7 : 0]     din56,
    input  [7 : 0]     din57,
    input  [7 : 0]     din58,
    input  [7 : 0]     din59,
    input  [7 : 0]     din60,
    input  [7 : 0]     din61,
    input  [7 : 0]     din62,
    input  [7 : 0]     din63,
    input  [7 : 0]     din64,
    input  [7 : 0]     din65,
    input  [7 : 0]     din66,
    input  [7 : 0]     din67,
    input  [7 : 0]     din68,
    input  [7 : 0]     din69,
    input  [7 : 0]     din70,
    input  [7 : 0]     din71,
    input  [7 : 0]     din72,
    input  [7 : 0]     din73,
    input  [7 : 0]     din74,
    input  [7 : 0]     din75,
    input  [7 : 0]     din76,
    input  [7 : 0]     din77,
    input  [7 : 0]     din78,
    input  [7 : 0]     din79,
    input  [7 : 0]     din80,
    input  [7 : 0]     din81,
    input  [7 : 0]     din82,
    input  [7 : 0]     din83,
    input  [7 : 0]     din84,
    input  [7 : 0]     din85,
    input  [7 : 0]     din86,
    input  [7 : 0]     din87,
    input  [7 : 0]     din88,
    input  [7 : 0]     din89,
    input  [7 : 0]     din90,
    input  [7 : 0]     din91,
    input  [7 : 0]     din92,
    input  [7 : 0]     din93,
    input  [7 : 0]     din94,
    input  [7 : 0]     din95,
    input  [7 : 0]     din96,
    input  [7 : 0]     din97,
    input  [7 : 0]     din98,
    input  [7 : 0]     din99,
    input  [7 : 0]     din100,
    input  [7 : 0]     din101,
    input  [7 : 0]     din102,
    input  [7 : 0]     din103,
    input  [7 : 0]     din104,
    input  [7 : 0]     din105,
    input  [7 : 0]     din106,
    input  [7 : 0]     din107,
    input  [7 : 0]     din108,
    input  [7 : 0]     din109,
    input  [7 : 0]     din110,
    input  [7 : 0]     din111,
    input  [7 : 0]     din112,
    input  [7 : 0]     din113,
    input  [7 : 0]     din114,
    input  [7 : 0]     din115,
    input  [7 : 0]     din116,
    input  [7 : 0]     din117,
    input  [7 : 0]     din118,
    input  [7 : 0]     din119,
    input  [7 : 0]     din120,
    input  [7 : 0]     din121,
    input  [7 : 0]     din122,
    input  [7 : 0]     din123,
    input  [7 : 0]     din124,
    input  [7 : 0]     din125,
    input  [7 : 0]     din126,
    input  [7 : 0]     din127,
    input  [7 : 0]     din128,
    input  [7 : 0]     din129,
    input  [7 : 0]     din130,
    input  [7 : 0]     din131,
    input  [7 : 0]     din132,
    input  [7 : 0]     din133,
    input  [7 : 0]     din134,
    input  [7 : 0]     din135,
    input  [7 : 0]     din136,
    input  [7 : 0]     din137,
    input  [7 : 0]     din138,
    input  [7 : 0]     din139,
    input  [7 : 0]     din140,
    input  [7 : 0]     din141,
    input  [7 : 0]     din142,
    input  [7 : 0]     din143,
    input  [7 : 0]     din144,
    input  [7 : 0]     din145,
    input  [7 : 0]     din146,
    input  [7 : 0]     din147,
    input  [7 : 0]     din148,
    input  [7 : 0]     din149,
    input  [7 : 0]     din150,
    input  [7 : 0]     din151,
    input  [7 : 0]     din152,
    input  [7 : 0]     din153,
    input  [7 : 0]     din154,
    input  [7 : 0]     din155,
    input  [7 : 0]     din156,
    input  [7 : 0]     din157,
    input  [7 : 0]     din158,
    input  [7 : 0]     din159,
    input  [7 : 0]     din160,
    input  [7 : 0]     din161,
    input  [7 : 0]     din162,
    input  [7 : 0]     din163,
    input  [7 : 0]     din164,
    input  [7 : 0]     din165,
    input  [7 : 0]     din166,
    input  [7 : 0]     din167,
    input  [7 : 0]     din168,
    input  [7 : 0]     din169,
    input  [7 : 0]     din170,
    input  [7 : 0]     din171,
    input  [7 : 0]     din172,
    input  [7 : 0]     din173,
    input  [7 : 0]     din174,
    input  [7 : 0]     din175,
    input  [7 : 0]     din176,
    input  [7 : 0]     din177,
    input  [7 : 0]     din178,
    input  [7 : 0]     din179,
    input  [7 : 0]     din180,
    input  [7 : 0]     din181,
    input  [7 : 0]     din182,
    input  [7 : 0]     din183,
    input  [7 : 0]     din184,
    input  [7 : 0]     din185,
    input  [7 : 0]     din186,
    input  [7 : 0]     din187,
    input  [7 : 0]     din188,
    input  [7 : 0]     din189,
    input  [7 : 0]     din190,
    input  [7 : 0]     din191,
    input  [7 : 0]     din192,
    input  [7 : 0]     din193,
    input  [7 : 0]     din194,
    input  [7 : 0]     din195,
    input  [7 : 0]     din196,
    input  [7 : 0]     din197,
    input  [7 : 0]     din198,
    input  [7 : 0]     din199,
    input  [7 : 0]     din200,
    input  [7 : 0]     din201,
    input  [7 : 0]     din202,
    input  [7 : 0]     din203,
    input  [7 : 0]     din204,
    input  [7 : 0]     din205,
    input  [7 : 0]     din206,
    input  [7 : 0]     din207,
    input  [7 : 0]     din208,
    input  [7 : 0]     din209,
    input  [7 : 0]     din210,
    input  [7 : 0]     din211,
    input  [7 : 0]     din212,
    input  [7 : 0]     din213,
    input  [7 : 0]     din214,
    input  [7 : 0]     din215,
    input  [7 : 0]     din216,
    input  [7 : 0]     din217,
    input  [7 : 0]     din218,
    input  [7 : 0]     din219,
    input  [7 : 0]     din220,
    input  [7 : 0]     din221,
    input  [7 : 0]     din222,
    input  [7 : 0]     din223,
    input  [7 : 0]     din224,
    input  [7 : 0]     din225,
    input  [7 : 0]     din226,
    input  [7 : 0]     din227,
    input  [7 : 0]     din228,
    input  [7 : 0]     din229,
    input  [7 : 0]     din230,
    input  [7 : 0]     din231,
    input  [7 : 0]     din232,
    input  [7 : 0]     din233,
    input  [7 : 0]     din234,
    input  [7 : 0]     din235,
    input  [7 : 0]     din236,
    input  [7 : 0]     din237,
    input  [7 : 0]     din238,
    input  [7 : 0]     din239,
    input  [7 : 0]     din240,
    input  [7 : 0]     din241,
    input  [7 : 0]     din242,
    input  [7 : 0]     din243,
    input  [7 : 0]     din244,
    input  [7 : 0]     din245,
    input  [7 : 0]     din246,
    input  [7 : 0]     din247,
    input  [7 : 0]     din248,
    input  [7 : 0]     din249,
    input  [7 : 0]     din250,
    input  [7 : 0]     din251,
    input  [7 : 0]     din252,
    input  [7 : 0]     din253,
    input  [7 : 0]     din254,
    input  [7 : 0]     din255,
    input  [7 : 0]    din256,
    output [7 : 0]   dout);

// puts internal signals
wire [7 : 0]     sel;
// level 1 signals
wire [7 : 0]         mux_1_0;
wire [7 : 0]         mux_1_1;
wire [7 : 0]         mux_1_2;
wire [7 : 0]         mux_1_3;
wire [7 : 0]         mux_1_4;
wire [7 : 0]         mux_1_5;
wire [7 : 0]         mux_1_6;
wire [7 : 0]         mux_1_7;
wire [7 : 0]         mux_1_8;
wire [7 : 0]         mux_1_9;
wire [7 : 0]         mux_1_10;
wire [7 : 0]         mux_1_11;
wire [7 : 0]         mux_1_12;
wire [7 : 0]         mux_1_13;
wire [7 : 0]         mux_1_14;
wire [7 : 0]         mux_1_15;
wire [7 : 0]         mux_1_16;
wire [7 : 0]         mux_1_17;
wire [7 : 0]         mux_1_18;
wire [7 : 0]         mux_1_19;
wire [7 : 0]         mux_1_20;
wire [7 : 0]         mux_1_21;
wire [7 : 0]         mux_1_22;
wire [7 : 0]         mux_1_23;
wire [7 : 0]         mux_1_24;
wire [7 : 0]         mux_1_25;
wire [7 : 0]         mux_1_26;
wire [7 : 0]         mux_1_27;
wire [7 : 0]         mux_1_28;
wire [7 : 0]         mux_1_29;
wire [7 : 0]         mux_1_30;
wire [7 : 0]         mux_1_31;
wire [7 : 0]         mux_1_32;
wire [7 : 0]         mux_1_33;
wire [7 : 0]         mux_1_34;
wire [7 : 0]         mux_1_35;
wire [7 : 0]         mux_1_36;
wire [7 : 0]         mux_1_37;
wire [7 : 0]         mux_1_38;
wire [7 : 0]         mux_1_39;
wire [7 : 0]         mux_1_40;
wire [7 : 0]         mux_1_41;
wire [7 : 0]         mux_1_42;
wire [7 : 0]         mux_1_43;
wire [7 : 0]         mux_1_44;
wire [7 : 0]         mux_1_45;
wire [7 : 0]         mux_1_46;
wire [7 : 0]         mux_1_47;
wire [7 : 0]         mux_1_48;
wire [7 : 0]         mux_1_49;
wire [7 : 0]         mux_1_50;
wire [7 : 0]         mux_1_51;
wire [7 : 0]         mux_1_52;
wire [7 : 0]         mux_1_53;
wire [7 : 0]         mux_1_54;
wire [7 : 0]         mux_1_55;
wire [7 : 0]         mux_1_56;
wire [7 : 0]         mux_1_57;
wire [7 : 0]         mux_1_58;
wire [7 : 0]         mux_1_59;
wire [7 : 0]         mux_1_60;
wire [7 : 0]         mux_1_61;
wire [7 : 0]         mux_1_62;
wire [7 : 0]         mux_1_63;
wire [7 : 0]         mux_1_64;
wire [7 : 0]         mux_1_65;
wire [7 : 0]         mux_1_66;
wire [7 : 0]         mux_1_67;
wire [7 : 0]         mux_1_68;
wire [7 : 0]         mux_1_69;
wire [7 : 0]         mux_1_70;
wire [7 : 0]         mux_1_71;
wire [7 : 0]         mux_1_72;
wire [7 : 0]         mux_1_73;
wire [7 : 0]         mux_1_74;
wire [7 : 0]         mux_1_75;
wire [7 : 0]         mux_1_76;
wire [7 : 0]         mux_1_77;
wire [7 : 0]         mux_1_78;
wire [7 : 0]         mux_1_79;
wire [7 : 0]         mux_1_80;
wire [7 : 0]         mux_1_81;
wire [7 : 0]         mux_1_82;
wire [7 : 0]         mux_1_83;
wire [7 : 0]         mux_1_84;
wire [7 : 0]         mux_1_85;
wire [7 : 0]         mux_1_86;
wire [7 : 0]         mux_1_87;
wire [7 : 0]         mux_1_88;
wire [7 : 0]         mux_1_89;
wire [7 : 0]         mux_1_90;
wire [7 : 0]         mux_1_91;
wire [7 : 0]         mux_1_92;
wire [7 : 0]         mux_1_93;
wire [7 : 0]         mux_1_94;
wire [7 : 0]         mux_1_95;
wire [7 : 0]         mux_1_96;
wire [7 : 0]         mux_1_97;
wire [7 : 0]         mux_1_98;
wire [7 : 0]         mux_1_99;
wire [7 : 0]         mux_1_100;
wire [7 : 0]         mux_1_101;
wire [7 : 0]         mux_1_102;
wire [7 : 0]         mux_1_103;
wire [7 : 0]         mux_1_104;
wire [7 : 0]         mux_1_105;
wire [7 : 0]         mux_1_106;
wire [7 : 0]         mux_1_107;
wire [7 : 0]         mux_1_108;
wire [7 : 0]         mux_1_109;
wire [7 : 0]         mux_1_110;
wire [7 : 0]         mux_1_111;
wire [7 : 0]         mux_1_112;
wire [7 : 0]         mux_1_113;
wire [7 : 0]         mux_1_114;
wire [7 : 0]         mux_1_115;
wire [7 : 0]         mux_1_116;
wire [7 : 0]         mux_1_117;
wire [7 : 0]         mux_1_118;
wire [7 : 0]         mux_1_119;
wire [7 : 0]         mux_1_120;
wire [7 : 0]         mux_1_121;
wire [7 : 0]         mux_1_122;
wire [7 : 0]         mux_1_123;
wire [7 : 0]         mux_1_124;
wire [7 : 0]         mux_1_125;
wire [7 : 0]         mux_1_126;
wire [7 : 0]         mux_1_127;
// level 2 signals
wire [7 : 0]         mux_2_0;
wire [7 : 0]         mux_2_1;
wire [7 : 0]         mux_2_2;
wire [7 : 0]         mux_2_3;
wire [7 : 0]         mux_2_4;
wire [7 : 0]         mux_2_5;
wire [7 : 0]         mux_2_6;
wire [7 : 0]         mux_2_7;
wire [7 : 0]         mux_2_8;
wire [7 : 0]         mux_2_9;
wire [7 : 0]         mux_2_10;
wire [7 : 0]         mux_2_11;
wire [7 : 0]         mux_2_12;
wire [7 : 0]         mux_2_13;
wire [7 : 0]         mux_2_14;
wire [7 : 0]         mux_2_15;
wire [7 : 0]         mux_2_16;
wire [7 : 0]         mux_2_17;
wire [7 : 0]         mux_2_18;
wire [7 : 0]         mux_2_19;
wire [7 : 0]         mux_2_20;
wire [7 : 0]         mux_2_21;
wire [7 : 0]         mux_2_22;
wire [7 : 0]         mux_2_23;
wire [7 : 0]         mux_2_24;
wire [7 : 0]         mux_2_25;
wire [7 : 0]         mux_2_26;
wire [7 : 0]         mux_2_27;
wire [7 : 0]         mux_2_28;
wire [7 : 0]         mux_2_29;
wire [7 : 0]         mux_2_30;
wire [7 : 0]         mux_2_31;
wire [7 : 0]         mux_2_32;
wire [7 : 0]         mux_2_33;
wire [7 : 0]         mux_2_34;
wire [7 : 0]         mux_2_35;
wire [7 : 0]         mux_2_36;
wire [7 : 0]         mux_2_37;
wire [7 : 0]         mux_2_38;
wire [7 : 0]         mux_2_39;
wire [7 : 0]         mux_2_40;
wire [7 : 0]         mux_2_41;
wire [7 : 0]         mux_2_42;
wire [7 : 0]         mux_2_43;
wire [7 : 0]         mux_2_44;
wire [7 : 0]         mux_2_45;
wire [7 : 0]         mux_2_46;
wire [7 : 0]         mux_2_47;
wire [7 : 0]         mux_2_48;
wire [7 : 0]         mux_2_49;
wire [7 : 0]         mux_2_50;
wire [7 : 0]         mux_2_51;
wire [7 : 0]         mux_2_52;
wire [7 : 0]         mux_2_53;
wire [7 : 0]         mux_2_54;
wire [7 : 0]         mux_2_55;
wire [7 : 0]         mux_2_56;
wire [7 : 0]         mux_2_57;
wire [7 : 0]         mux_2_58;
wire [7 : 0]         mux_2_59;
wire [7 : 0]         mux_2_60;
wire [7 : 0]         mux_2_61;
wire [7 : 0]         mux_2_62;
wire [7 : 0]         mux_2_63;
// level 3 signals
wire [7 : 0]         mux_3_0;
wire [7 : 0]         mux_3_1;
wire [7 : 0]         mux_3_2;
wire [7 : 0]         mux_3_3;
wire [7 : 0]         mux_3_4;
wire [7 : 0]         mux_3_5;
wire [7 : 0]         mux_3_6;
wire [7 : 0]         mux_3_7;
wire [7 : 0]         mux_3_8;
wire [7 : 0]         mux_3_9;
wire [7 : 0]         mux_3_10;
wire [7 : 0]         mux_3_11;
wire [7 : 0]         mux_3_12;
wire [7 : 0]         mux_3_13;
wire [7 : 0]         mux_3_14;
wire [7 : 0]         mux_3_15;
wire [7 : 0]         mux_3_16;
wire [7 : 0]         mux_3_17;
wire [7 : 0]         mux_3_18;
wire [7 : 0]         mux_3_19;
wire [7 : 0]         mux_3_20;
wire [7 : 0]         mux_3_21;
wire [7 : 0]         mux_3_22;
wire [7 : 0]         mux_3_23;
wire [7 : 0]         mux_3_24;
wire [7 : 0]         mux_3_25;
wire [7 : 0]         mux_3_26;
wire [7 : 0]         mux_3_27;
wire [7 : 0]         mux_3_28;
wire [7 : 0]         mux_3_29;
wire [7 : 0]         mux_3_30;
wire [7 : 0]         mux_3_31;
// level 4 signals
wire [7 : 0]         mux_4_0;
wire [7 : 0]         mux_4_1;
wire [7 : 0]         mux_4_2;
wire [7 : 0]         mux_4_3;
wire [7 : 0]         mux_4_4;
wire [7 : 0]         mux_4_5;
wire [7 : 0]         mux_4_6;
wire [7 : 0]         mux_4_7;
wire [7 : 0]         mux_4_8;
wire [7 : 0]         mux_4_9;
wire [7 : 0]         mux_4_10;
wire [7 : 0]         mux_4_11;
wire [7 : 0]         mux_4_12;
wire [7 : 0]         mux_4_13;
wire [7 : 0]         mux_4_14;
wire [7 : 0]         mux_4_15;
// level 5 signals
wire [7 : 0]         mux_5_0;
wire [7 : 0]         mux_5_1;
wire [7 : 0]         mux_5_2;
wire [7 : 0]         mux_5_3;
wire [7 : 0]         mux_5_4;
wire [7 : 0]         mux_5_5;
wire [7 : 0]         mux_5_6;
wire [7 : 0]         mux_5_7;
// level 6 signals
wire [7 : 0]         mux_6_0;
wire [7 : 0]         mux_6_1;
wire [7 : 0]         mux_6_2;
wire [7 : 0]         mux_6_3;
// level 7 signals
wire [7 : 0]         mux_7_0;
wire [7 : 0]         mux_7_1;
// level 8 signals
wire [7 : 0]         mux_8_0;

assign sel = din256;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;
assign mux_1_2 = (sel[0] == 0)? din4 : din5;
assign mux_1_3 = (sel[0] == 0)? din6 : din7;
assign mux_1_4 = (sel[0] == 0)? din8 : din9;
assign mux_1_5 = (sel[0] == 0)? din10 : din11;
assign mux_1_6 = (sel[0] == 0)? din12 : din13;
assign mux_1_7 = (sel[0] == 0)? din14 : din15;
assign mux_1_8 = (sel[0] == 0)? din16 : din17;
assign mux_1_9 = (sel[0] == 0)? din18 : din19;
assign mux_1_10 = (sel[0] == 0)? din20 : din21;
assign mux_1_11 = (sel[0] == 0)? din22 : din23;
assign mux_1_12 = (sel[0] == 0)? din24 : din25;
assign mux_1_13 = (sel[0] == 0)? din26 : din27;
assign mux_1_14 = (sel[0] == 0)? din28 : din29;
assign mux_1_15 = (sel[0] == 0)? din30 : din31;
assign mux_1_16 = (sel[0] == 0)? din32 : din33;
assign mux_1_17 = (sel[0] == 0)? din34 : din35;
assign mux_1_18 = (sel[0] == 0)? din36 : din37;
assign mux_1_19 = (sel[0] == 0)? din38 : din39;
assign mux_1_20 = (sel[0] == 0)? din40 : din41;
assign mux_1_21 = (sel[0] == 0)? din42 : din43;
assign mux_1_22 = (sel[0] == 0)? din44 : din45;
assign mux_1_23 = (sel[0] == 0)? din46 : din47;
assign mux_1_24 = (sel[0] == 0)? din48 : din49;
assign mux_1_25 = (sel[0] == 0)? din50 : din51;
assign mux_1_26 = (sel[0] == 0)? din52 : din53;
assign mux_1_27 = (sel[0] == 0)? din54 : din55;
assign mux_1_28 = (sel[0] == 0)? din56 : din57;
assign mux_1_29 = (sel[0] == 0)? din58 : din59;
assign mux_1_30 = (sel[0] == 0)? din60 : din61;
assign mux_1_31 = (sel[0] == 0)? din62 : din63;
assign mux_1_32 = (sel[0] == 0)? din64 : din65;
assign mux_1_33 = (sel[0] == 0)? din66 : din67;
assign mux_1_34 = (sel[0] == 0)? din68 : din69;
assign mux_1_35 = (sel[0] == 0)? din70 : din71;
assign mux_1_36 = (sel[0] == 0)? din72 : din73;
assign mux_1_37 = (sel[0] == 0)? din74 : din75;
assign mux_1_38 = (sel[0] == 0)? din76 : din77;
assign mux_1_39 = (sel[0] == 0)? din78 : din79;
assign mux_1_40 = (sel[0] == 0)? din80 : din81;
assign mux_1_41 = (sel[0] == 0)? din82 : din83;
assign mux_1_42 = (sel[0] == 0)? din84 : din85;
assign mux_1_43 = (sel[0] == 0)? din86 : din87;
assign mux_1_44 = (sel[0] == 0)? din88 : din89;
assign mux_1_45 = (sel[0] == 0)? din90 : din91;
assign mux_1_46 = (sel[0] == 0)? din92 : din93;
assign mux_1_47 = (sel[0] == 0)? din94 : din95;
assign mux_1_48 = (sel[0] == 0)? din96 : din97;
assign mux_1_49 = (sel[0] == 0)? din98 : din99;
assign mux_1_50 = (sel[0] == 0)? din100 : din101;
assign mux_1_51 = (sel[0] == 0)? din102 : din103;
assign mux_1_52 = (sel[0] == 0)? din104 : din105;
assign mux_1_53 = (sel[0] == 0)? din106 : din107;
assign mux_1_54 = (sel[0] == 0)? din108 : din109;
assign mux_1_55 = (sel[0] == 0)? din110 : din111;
assign mux_1_56 = (sel[0] == 0)? din112 : din113;
assign mux_1_57 = (sel[0] == 0)? din114 : din115;
assign mux_1_58 = (sel[0] == 0)? din116 : din117;
assign mux_1_59 = (sel[0] == 0)? din118 : din119;
assign mux_1_60 = (sel[0] == 0)? din120 : din121;
assign mux_1_61 = (sel[0] == 0)? din122 : din123;
assign mux_1_62 = (sel[0] == 0)? din124 : din125;
assign mux_1_63 = (sel[0] == 0)? din126 : din127;
assign mux_1_64 = (sel[0] == 0)? din128 : din129;
assign mux_1_65 = (sel[0] == 0)? din130 : din131;
assign mux_1_66 = (sel[0] == 0)? din132 : din133;
assign mux_1_67 = (sel[0] == 0)? din134 : din135;
assign mux_1_68 = (sel[0] == 0)? din136 : din137;
assign mux_1_69 = (sel[0] == 0)? din138 : din139;
assign mux_1_70 = (sel[0] == 0)? din140 : din141;
assign mux_1_71 = (sel[0] == 0)? din142 : din143;
assign mux_1_72 = (sel[0] == 0)? din144 : din145;
assign mux_1_73 = (sel[0] == 0)? din146 : din147;
assign mux_1_74 = (sel[0] == 0)? din148 : din149;
assign mux_1_75 = (sel[0] == 0)? din150 : din151;
assign mux_1_76 = (sel[0] == 0)? din152 : din153;
assign mux_1_77 = (sel[0] == 0)? din154 : din155;
assign mux_1_78 = (sel[0] == 0)? din156 : din157;
assign mux_1_79 = (sel[0] == 0)? din158 : din159;
assign mux_1_80 = (sel[0] == 0)? din160 : din161;
assign mux_1_81 = (sel[0] == 0)? din162 : din163;
assign mux_1_82 = (sel[0] == 0)? din164 : din165;
assign mux_1_83 = (sel[0] == 0)? din166 : din167;
assign mux_1_84 = (sel[0] == 0)? din168 : din169;
assign mux_1_85 = (sel[0] == 0)? din170 : din171;
assign mux_1_86 = (sel[0] == 0)? din172 : din173;
assign mux_1_87 = (sel[0] == 0)? din174 : din175;
assign mux_1_88 = (sel[0] == 0)? din176 : din177;
assign mux_1_89 = (sel[0] == 0)? din178 : din179;
assign mux_1_90 = (sel[0] == 0)? din180 : din181;
assign mux_1_91 = (sel[0] == 0)? din182 : din183;
assign mux_1_92 = (sel[0] == 0)? din184 : din185;
assign mux_1_93 = (sel[0] == 0)? din186 : din187;
assign mux_1_94 = (sel[0] == 0)? din188 : din189;
assign mux_1_95 = (sel[0] == 0)? din190 : din191;
assign mux_1_96 = (sel[0] == 0)? din192 : din193;
assign mux_1_97 = (sel[0] == 0)? din194 : din195;
assign mux_1_98 = (sel[0] == 0)? din196 : din197;
assign mux_1_99 = (sel[0] == 0)? din198 : din199;
assign mux_1_100 = (sel[0] == 0)? din200 : din201;
assign mux_1_101 = (sel[0] == 0)? din202 : din203;
assign mux_1_102 = (sel[0] == 0)? din204 : din205;
assign mux_1_103 = (sel[0] == 0)? din206 : din207;
assign mux_1_104 = (sel[0] == 0)? din208 : din209;
assign mux_1_105 = (sel[0] == 0)? din210 : din211;
assign mux_1_106 = (sel[0] == 0)? din212 : din213;
assign mux_1_107 = (sel[0] == 0)? din214 : din215;
assign mux_1_108 = (sel[0] == 0)? din216 : din217;
assign mux_1_109 = (sel[0] == 0)? din218 : din219;
assign mux_1_110 = (sel[0] == 0)? din220 : din221;
assign mux_1_111 = (sel[0] == 0)? din222 : din223;
assign mux_1_112 = (sel[0] == 0)? din224 : din225;
assign mux_1_113 = (sel[0] == 0)? din226 : din227;
assign mux_1_114 = (sel[0] == 0)? din228 : din229;
assign mux_1_115 = (sel[0] == 0)? din230 : din231;
assign mux_1_116 = (sel[0] == 0)? din232 : din233;
assign mux_1_117 = (sel[0] == 0)? din234 : din235;
assign mux_1_118 = (sel[0] == 0)? din236 : din237;
assign mux_1_119 = (sel[0] == 0)? din238 : din239;
assign mux_1_120 = (sel[0] == 0)? din240 : din241;
assign mux_1_121 = (sel[0] == 0)? din242 : din243;
assign mux_1_122 = (sel[0] == 0)? din244 : din245;
assign mux_1_123 = (sel[0] == 0)? din246 : din247;
assign mux_1_124 = (sel[0] == 0)? din248 : din249;
assign mux_1_125 = (sel[0] == 0)? din250 : din251;
assign mux_1_126 = (sel[0] == 0)? din252 : din253;
assign mux_1_127 = (sel[0] == 0)? din254 : din255;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;
assign mux_2_1 = (sel[1] == 0)? mux_1_2 : mux_1_3;
assign mux_2_2 = (sel[1] == 0)? mux_1_4 : mux_1_5;
assign mux_2_3 = (sel[1] == 0)? mux_1_6 : mux_1_7;
assign mux_2_4 = (sel[1] == 0)? mux_1_8 : mux_1_9;
assign mux_2_5 = (sel[1] == 0)? mux_1_10 : mux_1_11;
assign mux_2_6 = (sel[1] == 0)? mux_1_12 : mux_1_13;
assign mux_2_7 = (sel[1] == 0)? mux_1_14 : mux_1_15;
assign mux_2_8 = (sel[1] == 0)? mux_1_16 : mux_1_17;
assign mux_2_9 = (sel[1] == 0)? mux_1_18 : mux_1_19;
assign mux_2_10 = (sel[1] == 0)? mux_1_20 : mux_1_21;
assign mux_2_11 = (sel[1] == 0)? mux_1_22 : mux_1_23;
assign mux_2_12 = (sel[1] == 0)? mux_1_24 : mux_1_25;
assign mux_2_13 = (sel[1] == 0)? mux_1_26 : mux_1_27;
assign mux_2_14 = (sel[1] == 0)? mux_1_28 : mux_1_29;
assign mux_2_15 = (sel[1] == 0)? mux_1_30 : mux_1_31;
assign mux_2_16 = (sel[1] == 0)? mux_1_32 : mux_1_33;
assign mux_2_17 = (sel[1] == 0)? mux_1_34 : mux_1_35;
assign mux_2_18 = (sel[1] == 0)? mux_1_36 : mux_1_37;
assign mux_2_19 = (sel[1] == 0)? mux_1_38 : mux_1_39;
assign mux_2_20 = (sel[1] == 0)? mux_1_40 : mux_1_41;
assign mux_2_21 = (sel[1] == 0)? mux_1_42 : mux_1_43;
assign mux_2_22 = (sel[1] == 0)? mux_1_44 : mux_1_45;
assign mux_2_23 = (sel[1] == 0)? mux_1_46 : mux_1_47;
assign mux_2_24 = (sel[1] == 0)? mux_1_48 : mux_1_49;
assign mux_2_25 = (sel[1] == 0)? mux_1_50 : mux_1_51;
assign mux_2_26 = (sel[1] == 0)? mux_1_52 : mux_1_53;
assign mux_2_27 = (sel[1] == 0)? mux_1_54 : mux_1_55;
assign mux_2_28 = (sel[1] == 0)? mux_1_56 : mux_1_57;
assign mux_2_29 = (sel[1] == 0)? mux_1_58 : mux_1_59;
assign mux_2_30 = (sel[1] == 0)? mux_1_60 : mux_1_61;
assign mux_2_31 = (sel[1] == 0)? mux_1_62 : mux_1_63;
assign mux_2_32 = (sel[1] == 0)? mux_1_64 : mux_1_65;
assign mux_2_33 = (sel[1] == 0)? mux_1_66 : mux_1_67;
assign mux_2_34 = (sel[1] == 0)? mux_1_68 : mux_1_69;
assign mux_2_35 = (sel[1] == 0)? mux_1_70 : mux_1_71;
assign mux_2_36 = (sel[1] == 0)? mux_1_72 : mux_1_73;
assign mux_2_37 = (sel[1] == 0)? mux_1_74 : mux_1_75;
assign mux_2_38 = (sel[1] == 0)? mux_1_76 : mux_1_77;
assign mux_2_39 = (sel[1] == 0)? mux_1_78 : mux_1_79;
assign mux_2_40 = (sel[1] == 0)? mux_1_80 : mux_1_81;
assign mux_2_41 = (sel[1] == 0)? mux_1_82 : mux_1_83;
assign mux_2_42 = (sel[1] == 0)? mux_1_84 : mux_1_85;
assign mux_2_43 = (sel[1] == 0)? mux_1_86 : mux_1_87;
assign mux_2_44 = (sel[1] == 0)? mux_1_88 : mux_1_89;
assign mux_2_45 = (sel[1] == 0)? mux_1_90 : mux_1_91;
assign mux_2_46 = (sel[1] == 0)? mux_1_92 : mux_1_93;
assign mux_2_47 = (sel[1] == 0)? mux_1_94 : mux_1_95;
assign mux_2_48 = (sel[1] == 0)? mux_1_96 : mux_1_97;
assign mux_2_49 = (sel[1] == 0)? mux_1_98 : mux_1_99;
assign mux_2_50 = (sel[1] == 0)? mux_1_100 : mux_1_101;
assign mux_2_51 = (sel[1] == 0)? mux_1_102 : mux_1_103;
assign mux_2_52 = (sel[1] == 0)? mux_1_104 : mux_1_105;
assign mux_2_53 = (sel[1] == 0)? mux_1_106 : mux_1_107;
assign mux_2_54 = (sel[1] == 0)? mux_1_108 : mux_1_109;
assign mux_2_55 = (sel[1] == 0)? mux_1_110 : mux_1_111;
assign mux_2_56 = (sel[1] == 0)? mux_1_112 : mux_1_113;
assign mux_2_57 = (sel[1] == 0)? mux_1_114 : mux_1_115;
assign mux_2_58 = (sel[1] == 0)? mux_1_116 : mux_1_117;
assign mux_2_59 = (sel[1] == 0)? mux_1_118 : mux_1_119;
assign mux_2_60 = (sel[1] == 0)? mux_1_120 : mux_1_121;
assign mux_2_61 = (sel[1] == 0)? mux_1_122 : mux_1_123;
assign mux_2_62 = (sel[1] == 0)? mux_1_124 : mux_1_125;
assign mux_2_63 = (sel[1] == 0)? mux_1_126 : mux_1_127;

// Generate level 3 logic
assign mux_3_0 = (sel[2] == 0)? mux_2_0 : mux_2_1;
assign mux_3_1 = (sel[2] == 0)? mux_2_2 : mux_2_3;
assign mux_3_2 = (sel[2] == 0)? mux_2_4 : mux_2_5;
assign mux_3_3 = (sel[2] == 0)? mux_2_6 : mux_2_7;
assign mux_3_4 = (sel[2] == 0)? mux_2_8 : mux_2_9;
assign mux_3_5 = (sel[2] == 0)? mux_2_10 : mux_2_11;
assign mux_3_6 = (sel[2] == 0)? mux_2_12 : mux_2_13;
assign mux_3_7 = (sel[2] == 0)? mux_2_14 : mux_2_15;
assign mux_3_8 = (sel[2] == 0)? mux_2_16 : mux_2_17;
assign mux_3_9 = (sel[2] == 0)? mux_2_18 : mux_2_19;
assign mux_3_10 = (sel[2] == 0)? mux_2_20 : mux_2_21;
assign mux_3_11 = (sel[2] == 0)? mux_2_22 : mux_2_23;
assign mux_3_12 = (sel[2] == 0)? mux_2_24 : mux_2_25;
assign mux_3_13 = (sel[2] == 0)? mux_2_26 : mux_2_27;
assign mux_3_14 = (sel[2] == 0)? mux_2_28 : mux_2_29;
assign mux_3_15 = (sel[2] == 0)? mux_2_30 : mux_2_31;
assign mux_3_16 = (sel[2] == 0)? mux_2_32 : mux_2_33;
assign mux_3_17 = (sel[2] == 0)? mux_2_34 : mux_2_35;
assign mux_3_18 = (sel[2] == 0)? mux_2_36 : mux_2_37;
assign mux_3_19 = (sel[2] == 0)? mux_2_38 : mux_2_39;
assign mux_3_20 = (sel[2] == 0)? mux_2_40 : mux_2_41;
assign mux_3_21 = (sel[2] == 0)? mux_2_42 : mux_2_43;
assign mux_3_22 = (sel[2] == 0)? mux_2_44 : mux_2_45;
assign mux_3_23 = (sel[2] == 0)? mux_2_46 : mux_2_47;
assign mux_3_24 = (sel[2] == 0)? mux_2_48 : mux_2_49;
assign mux_3_25 = (sel[2] == 0)? mux_2_50 : mux_2_51;
assign mux_3_26 = (sel[2] == 0)? mux_2_52 : mux_2_53;
assign mux_3_27 = (sel[2] == 0)? mux_2_54 : mux_2_55;
assign mux_3_28 = (sel[2] == 0)? mux_2_56 : mux_2_57;
assign mux_3_29 = (sel[2] == 0)? mux_2_58 : mux_2_59;
assign mux_3_30 = (sel[2] == 0)? mux_2_60 : mux_2_61;
assign mux_3_31 = (sel[2] == 0)? mux_2_62 : mux_2_63;

// Generate level 4 logic
assign mux_4_0 = (sel[3] == 0)? mux_3_0 : mux_3_1;
assign mux_4_1 = (sel[3] == 0)? mux_3_2 : mux_3_3;
assign mux_4_2 = (sel[3] == 0)? mux_3_4 : mux_3_5;
assign mux_4_3 = (sel[3] == 0)? mux_3_6 : mux_3_7;
assign mux_4_4 = (sel[3] == 0)? mux_3_8 : mux_3_9;
assign mux_4_5 = (sel[3] == 0)? mux_3_10 : mux_3_11;
assign mux_4_6 = (sel[3] == 0)? mux_3_12 : mux_3_13;
assign mux_4_7 = (sel[3] == 0)? mux_3_14 : mux_3_15;
assign mux_4_8 = (sel[3] == 0)? mux_3_16 : mux_3_17;
assign mux_4_9 = (sel[3] == 0)? mux_3_18 : mux_3_19;
assign mux_4_10 = (sel[3] == 0)? mux_3_20 : mux_3_21;
assign mux_4_11 = (sel[3] == 0)? mux_3_22 : mux_3_23;
assign mux_4_12 = (sel[3] == 0)? mux_3_24 : mux_3_25;
assign mux_4_13 = (sel[3] == 0)? mux_3_26 : mux_3_27;
assign mux_4_14 = (sel[3] == 0)? mux_3_28 : mux_3_29;
assign mux_4_15 = (sel[3] == 0)? mux_3_30 : mux_3_31;

// Generate level 5 logic
assign mux_5_0 = (sel[4] == 0)? mux_4_0 : mux_4_1;
assign mux_5_1 = (sel[4] == 0)? mux_4_2 : mux_4_3;
assign mux_5_2 = (sel[4] == 0)? mux_4_4 : mux_4_5;
assign mux_5_3 = (sel[4] == 0)? mux_4_6 : mux_4_7;
assign mux_5_4 = (sel[4] == 0)? mux_4_8 : mux_4_9;
assign mux_5_5 = (sel[4] == 0)? mux_4_10 : mux_4_11;
assign mux_5_6 = (sel[4] == 0)? mux_4_12 : mux_4_13;
assign mux_5_7 = (sel[4] == 0)? mux_4_14 : mux_4_15;

// Generate level 6 logic
assign mux_6_0 = (sel[5] == 0)? mux_5_0 : mux_5_1;
assign mux_6_1 = (sel[5] == 0)? mux_5_2 : mux_5_3;
assign mux_6_2 = (sel[5] == 0)? mux_5_4 : mux_5_5;
assign mux_6_3 = (sel[5] == 0)? mux_5_6 : mux_5_7;

// Generate level 7 logic
assign mux_7_0 = (sel[6] == 0)? mux_6_0 : mux_6_1;
assign mux_7_1 = (sel[6] == 0)? mux_6_2 : mux_6_3;

// Generate level 8 logic
assign mux_8_0 = (sel[7] == 0)? mux_7_0 : mux_7_1;

// output logic
assign dout = mux_8_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/a3f1/hdl/verilog/ConvolutionInputGenerator_1_ConvolutionInputGbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module ConvolutionInputGenerator_1_ConvolutionInputGbkb_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 192;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];




always @(posedge clk)  
begin 
    if (ce0) begin
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module ConvolutionInputGenerator_1_ConvolutionInputGbkb(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd192;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



ConvolutionInputGenerator_1_ConvolutionInputGbkb_ram ConvolutionInputGenerator_1_ConvolutionInputGbkb_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_StreamingFCLayer_6jw.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

(* use_dsp = "no" *) module StreamingFCLayer_Batch_2_StreamingFCLayer_6jw_Mul_LUT_0(a, b, p);
input[8 - 1 : 0] a; 
input[4 - 1 : 0] b; 
output[12 - 1 : 0] p;

assign p = $signed(a) * $signed(b);
endmodule
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_StreamingFCLayer_6jw(
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



StreamingFCLayer_Batch_2_StreamingFCLayer_6jw_Mul_LUT_0 StreamingFCLayer_Batch_2_StreamingFCLayer_6jw_Mul_LUT_0_U(
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActXh4.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActXh4_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActXh4_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActXh4(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActXh4_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActXh4_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Activa.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module StreamingFCLayer_Batch_1_Matrix_Vector_Activa (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY,
        weight_V_V_TDATA,
        weight_V_V_TVALID,
        weight_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state6 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [15:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;
input  [63:0] weight_V_V_TDATA;
input   weight_V_V_TVALID;
output   weight_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;
reg weight_V_V_TREADY;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [5:0] threshs_m_thresholds_55_address0;
reg    threshs_m_thresholds_55_ce0;
wire   [15:0] threshs_m_thresholds_55_q0;
wire   [5:0] threshs_m_thresholds_54_address0;
reg    threshs_m_thresholds_54_ce0;
wire   [15:0] threshs_m_thresholds_54_q0;
wire   [5:0] threshs_m_thresholds_49_address0;
reg    threshs_m_thresholds_49_ce0;
wire   [15:0] threshs_m_thresholds_49_q0;
wire   [5:0] threshs_m_thresholds_48_address0;
reg    threshs_m_thresholds_48_ce0;
wire   [16:0] threshs_m_thresholds_48_q0;
wire   [5:0] threshs_m_thresholds_47_address0;
reg    threshs_m_thresholds_47_ce0;
wire   [16:0] threshs_m_thresholds_47_q0;
wire   [5:0] threshs_m_thresholds_46_address0;
reg    threshs_m_thresholds_46_ce0;
wire   [16:0] threshs_m_thresholds_46_q0;
wire   [5:0] threshs_m_thresholds_45_address0;
reg    threshs_m_thresholds_45_ce0;
wire   [16:0] threshs_m_thresholds_45_q0;
wire   [5:0] threshs_m_thresholds_44_address0;
reg    threshs_m_thresholds_44_ce0;
wire   [16:0] threshs_m_thresholds_44_q0;
wire   [5:0] threshs_m_thresholds_43_address0;
reg    threshs_m_thresholds_43_ce0;
wire   [16:0] threshs_m_thresholds_43_q0;
wire   [5:0] threshs_m_thresholds_42_address0;
reg    threshs_m_thresholds_42_ce0;
wire   [16:0] threshs_m_thresholds_42_q0;
wire   [5:0] threshs_m_thresholds_53_address0;
reg    threshs_m_thresholds_53_ce0;
wire   [16:0] threshs_m_thresholds_53_q0;
wire   [5:0] threshs_m_thresholds_52_address0;
reg    threshs_m_thresholds_52_ce0;
wire   [16:0] threshs_m_thresholds_52_q0;
wire   [5:0] threshs_m_thresholds_51_address0;
reg    threshs_m_thresholds_51_ce0;
wire   [16:0] threshs_m_thresholds_51_q0;
wire   [5:0] threshs_m_thresholds_50_address0;
reg    threshs_m_thresholds_50_ce0;
wire   [16:0] threshs_m_thresholds_50_q0;
wire   [5:0] threshs_m_thresholds_41_address0;
reg    threshs_m_thresholds_41_ce0;
wire   [17:0] threshs_m_thresholds_41_q0;
wire   [5:0] threshs_m_thresholds_40_address0;
reg    threshs_m_thresholds_40_ce0;
wire   [17:0] threshs_m_thresholds_40_q0;
wire   [5:0] threshs_m_thresholds_35_address0;
reg    threshs_m_thresholds_35_ce0;
wire   [17:0] threshs_m_thresholds_35_q0;
wire   [5:0] threshs_m_thresholds_34_address0;
reg    threshs_m_thresholds_34_ce0;
wire   [17:0] threshs_m_thresholds_34_q0;
wire   [5:0] threshs_m_thresholds_33_address0;
reg    threshs_m_thresholds_33_ce0;
wire   [17:0] threshs_m_thresholds_33_q0;
wire   [5:0] threshs_m_thresholds_32_address0;
reg    threshs_m_thresholds_32_ce0;
wire   [17:0] threshs_m_thresholds_32_q0;
wire   [5:0] threshs_m_thresholds_31_address0;
reg    threshs_m_thresholds_31_ce0;
wire   [17:0] threshs_m_thresholds_31_q0;
wire   [5:0] threshs_m_thresholds_30_address0;
reg    threshs_m_thresholds_30_ce0;
wire   [17:0] threshs_m_thresholds_30_q0;
wire   [5:0] threshs_m_thresholds_29_address0;
reg    threshs_m_thresholds_29_ce0;
wire   [17:0] threshs_m_thresholds_29_q0;
wire   [5:0] threshs_m_thresholds_28_address0;
reg    threshs_m_thresholds_28_ce0;
wire   [17:0] threshs_m_thresholds_28_q0;
wire   [5:0] threshs_m_thresholds_39_address0;
reg    threshs_m_thresholds_39_ce0;
wire   [17:0] threshs_m_thresholds_39_q0;
wire   [5:0] threshs_m_thresholds_38_address0;
reg    threshs_m_thresholds_38_ce0;
wire   [17:0] threshs_m_thresholds_38_q0;
wire   [5:0] threshs_m_thresholds_37_address0;
reg    threshs_m_thresholds_37_ce0;
wire   [17:0] threshs_m_thresholds_37_q0;
wire   [5:0] threshs_m_thresholds_36_address0;
reg    threshs_m_thresholds_36_ce0;
wire   [17:0] threshs_m_thresholds_36_q0;
wire   [5:0] threshs_m_thresholds_27_address0;
reg    threshs_m_thresholds_27_ce0;
wire   [16:0] threshs_m_thresholds_27_q0;
wire   [5:0] threshs_m_thresholds_26_address0;
reg    threshs_m_thresholds_26_ce0;
wire   [16:0] threshs_m_thresholds_26_q0;
wire   [5:0] threshs_m_thresholds_21_address0;
reg    threshs_m_thresholds_21_ce0;
wire   [16:0] threshs_m_thresholds_21_q0;
wire   [5:0] threshs_m_thresholds_20_address0;
reg    threshs_m_thresholds_20_ce0;
wire   [16:0] threshs_m_thresholds_20_q0;
wire   [5:0] threshs_m_thresholds_19_address0;
reg    threshs_m_thresholds_19_ce0;
wire   [16:0] threshs_m_thresholds_19_q0;
wire   [5:0] threshs_m_thresholds_18_address0;
reg    threshs_m_thresholds_18_ce0;
wire   [16:0] threshs_m_thresholds_18_q0;
wire   [5:0] threshs_m_thresholds_17_address0;
reg    threshs_m_thresholds_17_ce0;
wire   [16:0] threshs_m_thresholds_17_q0;
wire   [5:0] threshs_m_thresholds_16_address0;
reg    threshs_m_thresholds_16_ce0;
wire   [16:0] threshs_m_thresholds_16_q0;
wire   [5:0] threshs_m_thresholds_15_address0;
reg    threshs_m_thresholds_15_ce0;
wire   [15:0] threshs_m_thresholds_15_q0;
wire   [5:0] threshs_m_thresholds_14_address0;
reg    threshs_m_thresholds_14_ce0;
wire   [15:0] threshs_m_thresholds_14_q0;
wire   [5:0] threshs_m_thresholds_25_address0;
reg    threshs_m_thresholds_25_ce0;
wire   [16:0] threshs_m_thresholds_25_q0;
wire   [5:0] threshs_m_thresholds_24_address0;
reg    threshs_m_thresholds_24_ce0;
wire   [16:0] threshs_m_thresholds_24_q0;
wire   [5:0] threshs_m_thresholds_23_address0;
reg    threshs_m_thresholds_23_ce0;
wire   [16:0] threshs_m_thresholds_23_q0;
wire   [5:0] threshs_m_thresholds_22_address0;
reg    threshs_m_thresholds_22_ce0;
wire   [16:0] threshs_m_thresholds_22_q0;
wire   [5:0] threshs_m_thresholds_13_address0;
reg    threshs_m_thresholds_13_ce0;
wire   [17:0] threshs_m_thresholds_13_q0;
wire   [5:0] threshs_m_thresholds_12_address0;
reg    threshs_m_thresholds_12_ce0;
wire   [16:0] threshs_m_thresholds_12_q0;
wire   [5:0] threshs_m_thresholds_7_address0;
reg    threshs_m_thresholds_7_ce0;
wire   [16:0] threshs_m_thresholds_7_q0;
wire   [5:0] threshs_m_thresholds_6_address0;
reg    threshs_m_thresholds_6_ce0;
wire   [16:0] threshs_m_thresholds_6_q0;
wire   [5:0] threshs_m_thresholds_5_address0;
reg    threshs_m_thresholds_5_ce0;
wire   [16:0] threshs_m_thresholds_5_q0;
wire   [5:0] threshs_m_thresholds_4_address0;
reg    threshs_m_thresholds_4_ce0;
wire   [16:0] threshs_m_thresholds_4_q0;
wire   [5:0] threshs_m_thresholds_3_address0;
reg    threshs_m_thresholds_3_ce0;
wire   [16:0] threshs_m_thresholds_3_q0;
wire   [5:0] threshs_m_thresholds_2_address0;
reg    threshs_m_thresholds_2_ce0;
wire   [16:0] threshs_m_thresholds_2_q0;
wire   [5:0] threshs_m_thresholds_1_address0;
reg    threshs_m_thresholds_1_ce0;
wire   [16:0] threshs_m_thresholds_1_q0;
wire   [5:0] threshs_m_thresholds_address0;
reg    threshs_m_thresholds_ce0;
wire   [16:0] threshs_m_thresholds_q0;
wire   [5:0] threshs_m_thresholds_11_address0;
reg    threshs_m_thresholds_11_ce0;
wire   [16:0] threshs_m_thresholds_11_q0;
wire   [5:0] threshs_m_thresholds_10_address0;
reg    threshs_m_thresholds_10_ce0;
wire   [16:0] threshs_m_thresholds_10_q0;
wire   [5:0] threshs_m_thresholds_9_address0;
reg    threshs_m_thresholds_9_ce0;
wire   [17:0] threshs_m_thresholds_9_q0;
wire   [5:0] threshs_m_thresholds_8_address0;
reg    threshs_m_thresholds_8_ce0;
wire   [17:0] threshs_m_thresholds_8_q0;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln248_fu_5645_p2;
wire   [0:0] icmp_ln252_fu_5660_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter3;
reg   [0:0] icmp_ln289_reg_17768;
reg   [0:0] icmp_ln289_reg_17768_pp0_iter2_reg;
reg    weight_V_V_TDATA_blk_n;
reg   [15:0] i_0_reg_4465;
reg    ap_predicate_op1185_read_state2;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
reg    ap_block_state5_io;
reg    ap_block_pp0_stage0_11001;
wire   [15:0] i_fu_5651_p2;
wire   [15:0] inElem_V_1_fu_7401_p578;
wire   [9:0] trunc_ln321_fu_8559_p1;
wire   [0:0] icmp_ln271_fu_11446_p2;
reg   [0:0] icmp_ln271_reg_17680;
reg   [0:0] icmp_ln271_reg_17680_pp0_iter1_reg;
wire   [3:0] trunc_ln647_fu_11452_p1;
reg  signed [3:0] trunc_ln647_reg_17688;
reg  signed [3:0] p_Result_1_0_1_reg_17693;
reg  signed [3:0] p_Result_1_0_2_reg_17698;
reg  signed [3:0] p_Result_1_0_3_reg_17703;
reg  signed [3:0] p_Result_1_1_reg_17708;
reg  signed [3:0] p_Result_1_1_1_reg_17713;
reg  signed [3:0] p_Result_1_1_2_reg_17718;
reg  signed [3:0] p_Result_1_1_3_reg_17723;
reg  signed [3:0] p_Result_1_2_reg_17728;
reg  signed [3:0] p_Result_1_2_1_reg_17733;
reg  signed [3:0] p_Result_1_2_2_reg_17738;
reg  signed [3:0] p_Result_1_2_3_reg_17743;
reg  signed [3:0] p_Result_1_3_reg_17748;
reg  signed [3:0] p_Result_1_3_1_reg_17753;
reg  signed [3:0] p_Result_1_3_2_reg_17758;
reg  signed [3:0] p_Result_1_3_3_reg_17763;
wire   [0:0] icmp_ln289_fu_11612_p2;
reg   [0:0] icmp_ln289_reg_17768_pp0_iter1_reg;
wire  signed [7:0] mul_ln1352_1_fu_11661_p2;
reg  signed [7:0] mul_ln1352_1_reg_17772;
wire   [8:0] add_ln700_2_fu_11727_p2;
reg   [8:0] add_ln700_2_reg_17777;
wire  signed [7:0] mul_ln1352_5_fu_11749_p2;
reg  signed [7:0] mul_ln1352_5_reg_17782;
wire   [8:0] add_ln700_6_fu_11787_p2;
reg   [8:0] add_ln700_6_reg_17787;
wire  signed [7:0] mul_ln1352_9_fu_11809_p2;
reg  signed [7:0] mul_ln1352_9_reg_17792;
wire   [8:0] add_ln700_10_fu_11847_p2;
reg   [8:0] add_ln700_10_reg_17797;
wire  signed [7:0] mul_ln1352_13_fu_11869_p2;
reg  signed [7:0] mul_ln1352_13_reg_17802;
wire   [8:0] add_ln700_14_fu_11907_p2;
reg   [8:0] add_ln700_14_reg_17807;
wire   [0:0] icmp_ln899_fu_12137_p2;
reg   [0:0] icmp_ln899_reg_18092;
wire   [0:0] icmp_ln899_1_fu_12147_p2;
reg   [0:0] icmp_ln899_1_reg_18097;
wire   [0:0] icmp_ln899_2_fu_12157_p2;
reg   [0:0] icmp_ln899_2_reg_18102;
wire   [0:0] icmp_ln899_3_fu_12167_p2;
reg   [0:0] icmp_ln899_3_reg_18107;
wire   [0:0] icmp_ln899_4_fu_12177_p2;
reg   [0:0] icmp_ln899_4_reg_18112;
wire   [0:0] icmp_ln899_5_fu_12187_p2;
reg   [0:0] icmp_ln899_5_reg_18117;
wire   [0:0] icmp_ln899_6_fu_12197_p2;
reg   [0:0] icmp_ln899_6_reg_18122;
wire   [0:0] icmp_ln899_7_fu_12207_p2;
reg   [0:0] icmp_ln899_7_reg_18127;
wire   [0:0] icmp_ln899_8_fu_12217_p2;
reg   [0:0] icmp_ln899_8_reg_18132;
wire   [0:0] icmp_ln899_9_fu_12227_p2;
reg   [0:0] icmp_ln899_9_reg_18137;
wire   [0:0] icmp_ln899_10_fu_12237_p2;
reg   [0:0] icmp_ln899_10_reg_18142;
wire   [0:0] icmp_ln899_11_fu_12247_p2;
reg   [0:0] icmp_ln899_11_reg_18147;
wire   [0:0] icmp_ln899_12_fu_12257_p2;
reg   [0:0] icmp_ln899_12_reg_18152;
wire   [0:0] icmp_ln899_13_fu_12267_p2;
reg   [0:0] icmp_ln899_13_reg_18157;
wire   [0:0] icmp_ln899_14_fu_12273_p2;
reg   [0:0] icmp_ln899_14_reg_18162;
wire   [0:0] icmp_ln899_15_fu_12279_p2;
reg   [0:0] icmp_ln899_15_reg_18167;
wire   [0:0] icmp_ln899_16_fu_12285_p2;
reg   [0:0] icmp_ln899_16_reg_18172;
wire   [0:0] icmp_ln899_17_fu_12291_p2;
reg   [0:0] icmp_ln899_17_reg_18177;
wire   [0:0] icmp_ln899_18_fu_12297_p2;
reg   [0:0] icmp_ln899_18_reg_18182;
wire   [0:0] icmp_ln899_19_fu_12303_p2;
reg   [0:0] icmp_ln899_19_reg_18187;
wire   [0:0] icmp_ln899_20_fu_12309_p2;
reg   [0:0] icmp_ln899_20_reg_18192;
wire   [0:0] icmp_ln899_21_fu_12315_p2;
reg   [0:0] icmp_ln899_21_reg_18197;
wire   [0:0] icmp_ln899_22_fu_12321_p2;
reg   [0:0] icmp_ln899_22_reg_18202;
wire   [0:0] icmp_ln899_23_fu_12327_p2;
reg   [0:0] icmp_ln899_23_reg_18207;
wire   [0:0] icmp_ln899_24_fu_12333_p2;
reg   [0:0] icmp_ln899_24_reg_18212;
wire   [0:0] icmp_ln899_25_fu_12339_p2;
reg   [0:0] icmp_ln899_25_reg_18217;
wire   [0:0] icmp_ln899_26_fu_12345_p2;
reg   [0:0] icmp_ln899_26_reg_18222;
wire   [0:0] icmp_ln899_27_fu_12351_p2;
reg   [0:0] icmp_ln899_27_reg_18227;
wire   [0:0] icmp_ln899_28_fu_12361_p2;
reg   [0:0] icmp_ln899_28_reg_18232;
wire   [0:0] icmp_ln899_29_fu_12371_p2;
reg   [0:0] icmp_ln899_29_reg_18237;
wire   [0:0] icmp_ln899_30_fu_12381_p2;
reg   [0:0] icmp_ln899_30_reg_18242;
wire   [0:0] icmp_ln899_31_fu_12391_p2;
reg   [0:0] icmp_ln899_31_reg_18247;
wire   [0:0] icmp_ln899_32_fu_12401_p2;
reg   [0:0] icmp_ln899_32_reg_18252;
wire   [0:0] icmp_ln899_33_fu_12411_p2;
reg   [0:0] icmp_ln899_33_reg_18257;
wire   [0:0] icmp_ln899_34_fu_12421_p2;
reg   [0:0] icmp_ln899_34_reg_18262;
wire   [0:0] icmp_ln899_35_fu_12431_p2;
reg   [0:0] icmp_ln899_35_reg_18267;
wire   [0:0] icmp_ln899_36_fu_12441_p2;
reg   [0:0] icmp_ln899_36_reg_18272;
wire   [0:0] icmp_ln899_37_fu_12451_p2;
reg   [0:0] icmp_ln899_37_reg_18277;
wire   [0:0] icmp_ln899_38_fu_12461_p2;
reg   [0:0] icmp_ln899_38_reg_18282;
wire   [0:0] icmp_ln899_39_fu_12471_p2;
reg   [0:0] icmp_ln899_39_reg_18287;
wire   [0:0] icmp_ln899_40_fu_12481_p2;
reg   [0:0] icmp_ln899_40_reg_18292;
wire   [0:0] icmp_ln899_41_fu_12491_p2;
reg   [0:0] icmp_ln899_41_reg_18297;
wire   [0:0] icmp_ln899_42_fu_12497_p2;
reg   [0:0] icmp_ln899_42_reg_18302;
wire   [0:0] icmp_ln899_43_fu_12507_p2;
reg   [0:0] icmp_ln899_43_reg_18307;
wire   [0:0] icmp_ln899_44_fu_12517_p2;
reg   [0:0] icmp_ln899_44_reg_18312;
wire   [0:0] icmp_ln899_45_fu_12527_p2;
reg   [0:0] icmp_ln899_45_reg_18317;
wire   [0:0] icmp_ln899_46_fu_12537_p2;
reg   [0:0] icmp_ln899_46_reg_18322;
wire   [0:0] icmp_ln899_47_fu_12547_p2;
reg   [0:0] icmp_ln899_47_reg_18327;
wire   [0:0] icmp_ln899_48_fu_12557_p2;
reg   [0:0] icmp_ln899_48_reg_18332;
wire   [0:0] icmp_ln899_49_fu_12567_p2;
reg   [0:0] icmp_ln899_49_reg_18337;
wire   [0:0] icmp_ln899_50_fu_12577_p2;
reg   [0:0] icmp_ln899_50_reg_18342;
wire   [0:0] icmp_ln899_51_fu_12587_p2;
reg   [0:0] icmp_ln899_51_reg_18347;
wire   [0:0] icmp_ln899_52_fu_12597_p2;
reg   [0:0] icmp_ln899_52_reg_18352;
wire   [0:0] icmp_ln899_53_fu_12607_p2;
reg   [0:0] icmp_ln899_53_reg_18357;
wire   [0:0] icmp_ln899_54_fu_12613_p2;
reg   [0:0] icmp_ln899_54_reg_18362;
wire   [0:0] icmp_ln899_55_fu_12619_p2;
reg   [0:0] icmp_ln899_55_reg_18367;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
wire   [15:0] ap_phi_reg_pp0_iter0_act_m_val_V_reg_4476;
reg   [15:0] ap_phi_reg_pp0_iter1_act_m_val_V_reg_4476;
wire   [63:0] zext_ln142_fu_11916_p1;
reg   [17:0] accu_V_0_0_0_fu_1390;
wire   [17:0] accu_0_0_V_fu_12053_p2;
reg   [17:0] accu_V_0_1_0_fu_1394;
wire   [17:0] accu_0_1_V_fu_12071_p2;
reg   [17:0] accu_V_0_2_0_fu_1398;
wire   [17:0] accu_0_2_V_fu_12089_p2;
reg   [17:0] accu_V_0_3_0_fu_1402;
wire   [17:0] accu_0_3_V_fu_12107_p2;
reg   [31:0] sf_1_fu_1406;
wire   [31:0] sf_fu_11606_p2;
reg   [15:0] tmp_V_fu_1410;
reg   [15:0] tmp_V_1_fu_1414;
reg   [15:0] tmp_V_2_fu_1418;
reg   [15:0] tmp_V_4_fu_1422;
reg   [15:0] tmp_V_5_fu_1426;
reg   [15:0] tmp_V_6_fu_1430;
reg   [15:0] tmp_V_7_fu_1434;
reg   [15:0] tmp_V_8_fu_1438;
reg   [15:0] tmp_V_9_fu_1442;
reg   [15:0] tmp_V_10_fu_1446;
reg   [15:0] tmp_V_11_fu_1450;
reg   [15:0] tmp_V_12_fu_1454;
reg   [15:0] tmp_V_13_fu_1458;
reg   [15:0] tmp_V_14_fu_1462;
reg   [15:0] tmp_V_15_fu_1466;
reg   [15:0] tmp_V_16_fu_1470;
reg   [15:0] tmp_V_17_fu_1474;
reg   [15:0] tmp_V_18_fu_1478;
reg   [15:0] tmp_V_19_fu_1482;
reg   [15:0] tmp_V_20_fu_1486;
reg   [15:0] tmp_V_21_fu_1490;
reg   [15:0] tmp_V_22_fu_1494;
reg   [15:0] tmp_V_23_fu_1498;
reg   [15:0] tmp_V_24_fu_1502;
reg   [15:0] tmp_V_25_fu_1506;
reg   [15:0] tmp_V_26_fu_1510;
reg   [15:0] tmp_V_27_fu_1514;
reg   [15:0] tmp_V_28_fu_1518;
reg   [15:0] tmp_V_29_fu_1522;
reg   [15:0] tmp_V_30_fu_1526;
reg   [15:0] tmp_V_31_fu_1530;
reg   [15:0] tmp_V_32_fu_1534;
reg   [15:0] tmp_V_33_fu_1538;
reg   [15:0] tmp_V_34_fu_1542;
reg   [15:0] tmp_V_35_fu_1546;
reg   [15:0] tmp_V_36_fu_1550;
reg   [15:0] tmp_V_37_fu_1554;
reg   [15:0] tmp_V_38_fu_1558;
reg   [15:0] tmp_V_39_fu_1562;
reg   [15:0] tmp_V_40_fu_1566;
reg   [15:0] tmp_V_41_fu_1570;
reg   [15:0] tmp_V_42_fu_1574;
reg   [15:0] tmp_V_43_fu_1578;
reg   [15:0] tmp_V_44_fu_1582;
reg   [15:0] tmp_V_45_fu_1586;
reg   [15:0] tmp_V_46_fu_1590;
reg   [15:0] tmp_V_47_fu_1594;
reg   [15:0] tmp_V_48_fu_1598;
reg   [15:0] tmp_V_49_fu_1602;
reg   [15:0] tmp_V_50_fu_1606;
reg   [15:0] tmp_V_51_fu_1610;
reg   [15:0] tmp_V_52_fu_1614;
reg   [15:0] tmp_V_53_fu_1618;
reg   [15:0] tmp_V_54_fu_1622;
reg   [15:0] tmp_V_55_fu_1626;
reg   [15:0] tmp_V_56_fu_1630;
reg   [15:0] tmp_V_57_fu_1634;
reg   [15:0] tmp_V_58_fu_1638;
reg   [15:0] tmp_V_59_fu_1642;
reg   [15:0] tmp_V_60_fu_1646;
reg   [15:0] tmp_V_61_fu_1650;
reg   [15:0] tmp_V_62_fu_1654;
reg   [15:0] tmp_V_63_fu_1658;
reg   [15:0] tmp_V_64_fu_1662;
reg   [15:0] tmp_V_65_fu_1666;
reg   [15:0] tmp_V_66_fu_1670;
reg   [15:0] tmp_V_67_fu_1674;
reg   [15:0] tmp_V_68_fu_1678;
reg   [15:0] tmp_V_69_fu_1682;
reg   [15:0] tmp_V_70_fu_1686;
reg   [15:0] tmp_V_71_fu_1690;
reg   [15:0] tmp_V_72_fu_1694;
reg   [15:0] tmp_V_73_fu_1698;
reg   [15:0] tmp_V_74_fu_1702;
reg   [15:0] tmp_V_75_fu_1706;
reg   [15:0] tmp_V_76_fu_1710;
reg   [15:0] tmp_V_77_fu_1714;
reg   [15:0] tmp_V_78_fu_1718;
reg   [15:0] tmp_V_79_fu_1722;
reg   [15:0] tmp_V_80_fu_1726;
reg   [15:0] tmp_V_81_fu_1730;
reg   [15:0] tmp_V_82_fu_1734;
reg   [15:0] tmp_V_83_fu_1738;
reg   [15:0] tmp_V_84_fu_1742;
reg   [15:0] tmp_V_85_fu_1746;
reg   [15:0] tmp_V_86_fu_1750;
reg   [15:0] tmp_V_87_fu_1754;
reg   [15:0] tmp_V_88_fu_1758;
reg   [15:0] tmp_V_89_fu_1762;
reg   [15:0] tmp_V_90_fu_1766;
reg   [15:0] tmp_V_91_fu_1770;
reg   [15:0] tmp_V_92_fu_1774;
reg   [15:0] tmp_V_93_fu_1778;
reg   [15:0] tmp_V_94_fu_1782;
reg   [15:0] tmp_V_95_fu_1786;
reg   [15:0] tmp_V_96_fu_1790;
reg   [15:0] tmp_V_97_fu_1794;
reg   [15:0] tmp_V_98_fu_1798;
reg   [15:0] tmp_V_99_fu_1802;
reg   [15:0] tmp_V_100_fu_1806;
reg   [15:0] tmp_V_101_fu_1810;
reg   [15:0] tmp_V_102_fu_1814;
reg   [15:0] tmp_V_103_fu_1818;
reg   [15:0] tmp_V_104_fu_1822;
reg   [15:0] tmp_V_105_fu_1826;
reg   [15:0] tmp_V_106_fu_1830;
reg   [15:0] tmp_V_107_fu_1834;
reg   [15:0] tmp_V_108_fu_1838;
reg   [15:0] tmp_V_109_fu_1842;
reg   [15:0] tmp_V_110_fu_1846;
reg   [15:0] tmp_V_111_fu_1850;
reg   [15:0] tmp_V_112_fu_1854;
reg   [15:0] tmp_V_113_fu_1858;
reg   [15:0] tmp_V_114_fu_1862;
reg   [15:0] tmp_V_115_fu_1866;
reg   [15:0] tmp_V_116_fu_1870;
reg   [15:0] tmp_V_117_fu_1874;
reg   [15:0] tmp_V_118_fu_1878;
reg   [15:0] tmp_V_119_fu_1882;
reg   [15:0] tmp_V_120_fu_1886;
reg   [15:0] tmp_V_121_fu_1890;
reg   [15:0] tmp_V_122_fu_1894;
reg   [15:0] tmp_V_123_fu_1898;
reg   [15:0] tmp_V_124_fu_1902;
reg   [15:0] tmp_V_125_fu_1906;
reg   [15:0] tmp_V_126_fu_1910;
reg   [15:0] tmp_V_127_fu_1914;
reg   [15:0] tmp_V_128_fu_1918;
reg   [15:0] tmp_V_129_fu_1922;
reg   [15:0] tmp_V_130_fu_1926;
reg   [15:0] tmp_V_131_fu_1930;
reg   [15:0] tmp_V_132_fu_1934;
reg   [15:0] tmp_V_133_fu_1938;
reg   [15:0] tmp_V_134_fu_1942;
reg   [15:0] tmp_V_135_fu_1946;
reg   [15:0] tmp_V_136_fu_1950;
reg   [15:0] tmp_V_137_fu_1954;
reg   [15:0] tmp_V_138_fu_1958;
reg   [15:0] tmp_V_139_fu_1962;
reg   [15:0] tmp_V_140_fu_1966;
reg   [15:0] tmp_V_141_fu_1970;
reg   [15:0] tmp_V_142_fu_1974;
reg   [15:0] tmp_V_143_fu_1978;
reg   [15:0] tmp_V_144_fu_1982;
reg   [15:0] tmp_V_145_fu_1986;
reg   [15:0] tmp_V_146_fu_1990;
reg   [15:0] tmp_V_147_fu_1994;
reg   [15:0] tmp_V_148_fu_1998;
reg   [15:0] tmp_V_149_fu_2002;
reg   [15:0] tmp_V_150_fu_2006;
reg   [15:0] tmp_V_151_fu_2010;
reg   [15:0] tmp_V_152_fu_2014;
reg   [15:0] tmp_V_153_fu_2018;
reg   [15:0] tmp_V_154_fu_2022;
reg   [15:0] tmp_V_155_fu_2026;
reg   [15:0] tmp_V_156_fu_2030;
reg   [15:0] tmp_V_157_fu_2034;
reg   [15:0] tmp_V_158_fu_2038;
reg   [15:0] tmp_V_159_fu_2042;
reg   [15:0] tmp_V_160_fu_2046;
reg   [15:0] tmp_V_161_fu_2050;
reg   [15:0] tmp_V_162_fu_2054;
reg   [15:0] tmp_V_163_fu_2058;
reg   [15:0] tmp_V_164_fu_2062;
reg   [15:0] tmp_V_165_fu_2066;
reg   [15:0] tmp_V_166_fu_2070;
reg   [15:0] tmp_V_167_fu_2074;
reg   [15:0] tmp_V_168_fu_2078;
reg   [15:0] tmp_V_169_fu_2082;
reg   [15:0] tmp_V_170_fu_2086;
reg   [15:0] tmp_V_171_fu_2090;
reg   [15:0] tmp_V_172_fu_2094;
reg   [15:0] tmp_V_173_fu_2098;
reg   [15:0] tmp_V_174_fu_2102;
reg   [15:0] tmp_V_175_fu_2106;
reg   [15:0] tmp_V_176_fu_2110;
reg   [15:0] tmp_V_177_fu_2114;
reg   [15:0] tmp_V_178_fu_2118;
reg   [15:0] tmp_V_179_fu_2122;
reg   [15:0] tmp_V_180_fu_2126;
reg   [15:0] tmp_V_181_fu_2130;
reg   [15:0] tmp_V_182_fu_2134;
reg   [15:0] tmp_V_183_fu_2138;
reg   [15:0] tmp_V_184_fu_2142;
reg   [15:0] tmp_V_185_fu_2146;
reg   [15:0] tmp_V_186_fu_2150;
reg   [15:0] tmp_V_187_fu_2154;
reg   [15:0] tmp_V_188_fu_2158;
reg   [15:0] tmp_V_189_fu_2162;
reg   [15:0] tmp_V_190_fu_2166;
reg   [15:0] tmp_V_191_fu_2170;
reg   [15:0] tmp_V_192_fu_2174;
reg   [15:0] tmp_V_193_fu_2178;
reg   [15:0] tmp_V_194_fu_2182;
reg   [15:0] tmp_V_195_fu_2186;
reg   [15:0] tmp_V_196_fu_2190;
reg   [15:0] tmp_V_197_fu_2194;
reg   [15:0] tmp_V_198_fu_2198;
reg   [15:0] tmp_V_199_fu_2202;
reg   [15:0] tmp_V_200_fu_2206;
reg   [15:0] tmp_V_201_fu_2210;
reg   [15:0] tmp_V_202_fu_2214;
reg   [15:0] tmp_V_203_fu_2218;
reg   [15:0] tmp_V_204_fu_2222;
reg   [15:0] tmp_V_205_fu_2226;
reg   [15:0] tmp_V_206_fu_2230;
reg   [15:0] tmp_V_207_fu_2234;
reg   [15:0] tmp_V_208_fu_2238;
reg   [15:0] tmp_V_209_fu_2242;
reg   [15:0] tmp_V_210_fu_2246;
reg   [15:0] tmp_V_211_fu_2250;
reg   [15:0] tmp_V_212_fu_2254;
reg   [15:0] tmp_V_213_fu_2258;
reg   [15:0] tmp_V_214_fu_2262;
reg   [15:0] tmp_V_215_fu_2266;
reg   [15:0] tmp_V_216_fu_2270;
reg   [15:0] tmp_V_217_fu_2274;
reg   [15:0] tmp_V_218_fu_2278;
reg   [15:0] tmp_V_219_fu_2282;
reg   [15:0] tmp_V_220_fu_2286;
reg   [15:0] tmp_V_221_fu_2290;
reg   [15:0] tmp_V_222_fu_2294;
reg   [15:0] tmp_V_223_fu_2298;
reg   [15:0] tmp_V_224_fu_2302;
reg   [15:0] tmp_V_225_fu_2306;
reg   [15:0] tmp_V_226_fu_2310;
reg   [15:0] tmp_V_227_fu_2314;
reg   [15:0] tmp_V_228_fu_2318;
reg   [15:0] tmp_V_229_fu_2322;
reg   [15:0] tmp_V_230_fu_2326;
reg   [15:0] tmp_V_231_fu_2330;
reg   [15:0] tmp_V_232_fu_2334;
reg   [15:0] tmp_V_233_fu_2338;
reg   [15:0] tmp_V_234_fu_2342;
reg   [15:0] tmp_V_235_fu_2346;
reg   [15:0] tmp_V_236_fu_2350;
reg   [15:0] tmp_V_237_fu_2354;
reg   [15:0] tmp_V_238_fu_2358;
reg   [15:0] tmp_V_239_fu_2362;
reg   [15:0] tmp_V_240_fu_2366;
reg   [15:0] tmp_V_241_fu_2370;
reg   [15:0] tmp_V_242_fu_2374;
reg   [15:0] tmp_V_243_fu_2378;
reg   [15:0] tmp_V_244_fu_2382;
reg   [15:0] tmp_V_245_fu_2386;
reg   [15:0] tmp_V_246_fu_2390;
reg   [15:0] tmp_V_247_fu_2394;
reg   [15:0] tmp_V_248_fu_2398;
reg   [15:0] tmp_V_249_fu_2402;
reg   [15:0] tmp_V_250_fu_2406;
reg   [15:0] tmp_V_251_fu_2410;
reg   [15:0] tmp_V_252_fu_2414;
reg   [15:0] tmp_V_253_fu_2418;
reg   [15:0] tmp_V_254_fu_2422;
reg   [15:0] tmp_V_255_fu_2426;
reg   [15:0] tmp_V_256_fu_2430;
reg   [15:0] tmp_V_257_fu_2434;
reg   [15:0] tmp_V_258_fu_2438;
reg   [15:0] tmp_V_259_fu_2442;
reg   [15:0] tmp_V_260_fu_2446;
reg   [15:0] tmp_V_261_fu_2450;
reg   [15:0] tmp_V_262_fu_2454;
reg   [15:0] tmp_V_263_fu_2458;
reg   [15:0] tmp_V_264_fu_2462;
reg   [15:0] tmp_V_265_fu_2466;
reg   [15:0] tmp_V_266_fu_2470;
reg   [15:0] tmp_V_267_fu_2474;
reg   [15:0] tmp_V_268_fu_2478;
reg   [15:0] tmp_V_269_fu_2482;
reg   [15:0] tmp_V_270_fu_2486;
reg   [15:0] tmp_V_271_fu_2490;
reg   [15:0] tmp_V_272_fu_2494;
reg   [15:0] tmp_V_273_fu_2498;
reg   [15:0] tmp_V_274_fu_2502;
reg   [15:0] tmp_V_275_fu_2506;
reg   [15:0] tmp_V_276_fu_2510;
reg   [15:0] tmp_V_277_fu_2514;
reg   [15:0] tmp_V_278_fu_2518;
reg   [15:0] tmp_V_279_fu_2522;
reg   [15:0] tmp_V_280_fu_2526;
reg   [15:0] tmp_V_281_fu_2530;
reg   [15:0] tmp_V_282_fu_2534;
reg   [15:0] tmp_V_283_fu_2538;
reg   [15:0] tmp_V_284_fu_2542;
reg   [15:0] tmp_V_285_fu_2546;
reg   [15:0] tmp_V_286_fu_2550;
reg   [15:0] tmp_V_287_fu_2554;
reg   [15:0] tmp_V_288_fu_2558;
reg   [15:0] tmp_V_289_fu_2562;
reg   [15:0] tmp_V_290_fu_2566;
reg   [15:0] tmp_V_291_fu_2570;
reg   [15:0] tmp_V_292_fu_2574;
reg   [15:0] tmp_V_293_fu_2578;
reg   [15:0] tmp_V_294_fu_2582;
reg   [15:0] tmp_V_295_fu_2586;
reg   [15:0] tmp_V_296_fu_2590;
reg   [15:0] tmp_V_297_fu_2594;
reg   [15:0] tmp_V_298_fu_2598;
reg   [15:0] tmp_V_299_fu_2602;
reg   [15:0] tmp_V_300_fu_2606;
reg   [15:0] tmp_V_301_fu_2610;
reg   [15:0] tmp_V_302_fu_2614;
reg   [15:0] tmp_V_303_fu_2618;
reg   [15:0] tmp_V_304_fu_2622;
reg   [15:0] tmp_V_305_fu_2626;
reg   [15:0] tmp_V_306_fu_2630;
reg   [15:0] tmp_V_307_fu_2634;
reg   [15:0] tmp_V_308_fu_2638;
reg   [15:0] tmp_V_309_fu_2642;
reg   [15:0] tmp_V_310_fu_2646;
reg   [15:0] tmp_V_311_fu_2650;
reg   [15:0] tmp_V_312_fu_2654;
reg   [15:0] tmp_V_313_fu_2658;
reg   [15:0] tmp_V_314_fu_2662;
reg   [15:0] tmp_V_315_fu_2666;
reg   [15:0] tmp_V_316_fu_2670;
reg   [15:0] tmp_V_317_fu_2674;
reg   [15:0] tmp_V_318_fu_2678;
reg   [15:0] tmp_V_319_fu_2682;
reg   [15:0] tmp_V_320_fu_2686;
reg   [15:0] tmp_V_321_fu_2690;
reg   [15:0] tmp_V_322_fu_2694;
reg   [15:0] tmp_V_323_fu_2698;
reg   [15:0] tmp_V_324_fu_2702;
reg   [15:0] tmp_V_325_fu_2706;
reg   [15:0] tmp_V_326_fu_2710;
reg   [15:0] tmp_V_327_fu_2714;
reg   [15:0] tmp_V_328_fu_2718;
reg   [15:0] tmp_V_329_fu_2722;
reg   [15:0] tmp_V_330_fu_2726;
reg   [15:0] tmp_V_331_fu_2730;
reg   [15:0] tmp_V_332_fu_2734;
reg   [15:0] tmp_V_333_fu_2738;
reg   [15:0] tmp_V_334_fu_2742;
reg   [15:0] tmp_V_335_fu_2746;
reg   [15:0] tmp_V_336_fu_2750;
reg   [15:0] tmp_V_337_fu_2754;
reg   [15:0] tmp_V_338_fu_2758;
reg   [15:0] tmp_V_339_fu_2762;
reg   [15:0] tmp_V_340_fu_2766;
reg   [15:0] tmp_V_341_fu_2770;
reg   [15:0] tmp_V_342_fu_2774;
reg   [15:0] tmp_V_343_fu_2778;
reg   [15:0] tmp_V_344_fu_2782;
reg   [15:0] tmp_V_345_fu_2786;
reg   [15:0] tmp_V_346_fu_2790;
reg   [15:0] tmp_V_347_fu_2794;
reg   [15:0] tmp_V_348_fu_2798;
reg   [15:0] tmp_V_349_fu_2802;
reg   [15:0] tmp_V_350_fu_2806;
reg   [15:0] tmp_V_351_fu_2810;
reg   [15:0] tmp_V_352_fu_2814;
reg   [15:0] tmp_V_353_fu_2818;
reg   [15:0] tmp_V_354_fu_2822;
reg   [15:0] tmp_V_355_fu_2826;
reg   [15:0] tmp_V_356_fu_2830;
reg   [15:0] tmp_V_357_fu_2834;
reg   [15:0] tmp_V_358_fu_2838;
reg   [15:0] tmp_V_359_fu_2842;
reg   [15:0] tmp_V_360_fu_2846;
reg   [15:0] tmp_V_361_fu_2850;
reg   [15:0] tmp_V_362_fu_2854;
reg   [15:0] tmp_V_363_fu_2858;
reg   [15:0] tmp_V_364_fu_2862;
reg   [15:0] tmp_V_365_fu_2866;
reg   [15:0] tmp_V_366_fu_2870;
reg   [15:0] tmp_V_367_fu_2874;
reg   [15:0] tmp_V_368_fu_2878;
reg   [15:0] tmp_V_369_fu_2882;
reg   [15:0] tmp_V_370_fu_2886;
reg   [15:0] tmp_V_371_fu_2890;
reg   [15:0] tmp_V_372_fu_2894;
reg   [15:0] tmp_V_373_fu_2898;
reg   [15:0] tmp_V_374_fu_2902;
reg   [15:0] tmp_V_375_fu_2906;
reg   [15:0] tmp_V_376_fu_2910;
reg   [15:0] tmp_V_377_fu_2914;
reg   [15:0] tmp_V_378_fu_2918;
reg   [15:0] tmp_V_379_fu_2922;
reg   [15:0] tmp_V_380_fu_2926;
reg   [15:0] tmp_V_381_fu_2930;
reg   [15:0] tmp_V_382_fu_2934;
reg   [15:0] tmp_V_383_fu_2938;
reg   [15:0] tmp_V_384_fu_2942;
reg   [15:0] tmp_V_385_fu_2946;
reg   [15:0] tmp_V_386_fu_2950;
reg   [15:0] tmp_V_387_fu_2954;
reg   [15:0] tmp_V_388_fu_2958;
reg   [15:0] tmp_V_389_fu_2962;
reg   [15:0] tmp_V_390_fu_2966;
reg   [15:0] tmp_V_391_fu_2970;
reg   [15:0] tmp_V_392_fu_2974;
reg   [15:0] tmp_V_393_fu_2978;
reg   [15:0] tmp_V_394_fu_2982;
reg   [15:0] tmp_V_395_fu_2986;
reg   [15:0] tmp_V_396_fu_2990;
reg   [15:0] tmp_V_397_fu_2994;
reg   [15:0] tmp_V_398_fu_2998;
reg   [15:0] tmp_V_399_fu_3002;
reg   [15:0] tmp_V_400_fu_3006;
reg   [15:0] tmp_V_401_fu_3010;
reg   [15:0] tmp_V_402_fu_3014;
reg   [15:0] tmp_V_403_fu_3018;
reg   [15:0] tmp_V_404_fu_3022;
reg   [15:0] tmp_V_405_fu_3026;
reg   [15:0] tmp_V_406_fu_3030;
reg   [15:0] tmp_V_407_fu_3034;
reg   [15:0] tmp_V_408_fu_3038;
reg   [15:0] tmp_V_409_fu_3042;
reg   [15:0] tmp_V_410_fu_3046;
reg   [15:0] tmp_V_411_fu_3050;
reg   [15:0] tmp_V_412_fu_3054;
reg   [15:0] tmp_V_413_fu_3058;
reg   [15:0] tmp_V_414_fu_3062;
reg   [15:0] tmp_V_415_fu_3066;
reg   [15:0] tmp_V_416_fu_3070;
reg   [15:0] tmp_V_417_fu_3074;
reg   [15:0] tmp_V_418_fu_3078;
reg   [15:0] tmp_V_419_fu_3082;
reg   [15:0] tmp_V_420_fu_3086;
reg   [15:0] tmp_V_421_fu_3090;
reg   [15:0] tmp_V_422_fu_3094;
reg   [15:0] tmp_V_423_fu_3098;
reg   [15:0] tmp_V_424_fu_3102;
reg   [15:0] tmp_V_425_fu_3106;
reg   [15:0] tmp_V_426_fu_3110;
reg   [15:0] tmp_V_427_fu_3114;
reg   [15:0] tmp_V_428_fu_3118;
reg   [15:0] tmp_V_429_fu_3122;
reg   [15:0] tmp_V_430_fu_3126;
reg   [15:0] tmp_V_431_fu_3130;
reg   [15:0] tmp_V_432_fu_3134;
reg   [15:0] tmp_V_433_fu_3138;
reg   [15:0] tmp_V_434_fu_3142;
reg   [15:0] tmp_V_435_fu_3146;
reg   [15:0] tmp_V_436_fu_3150;
reg   [15:0] tmp_V_437_fu_3154;
reg   [15:0] tmp_V_438_fu_3158;
reg   [15:0] tmp_V_439_fu_3162;
reg   [15:0] tmp_V_440_fu_3166;
reg   [15:0] tmp_V_441_fu_3170;
reg   [15:0] tmp_V_442_fu_3174;
reg   [15:0] tmp_V_443_fu_3178;
reg   [15:0] tmp_V_444_fu_3182;
reg   [15:0] tmp_V_445_fu_3186;
reg   [15:0] tmp_V_446_fu_3190;
reg   [15:0] tmp_V_447_fu_3194;
reg   [15:0] tmp_V_448_fu_3198;
reg   [15:0] tmp_V_449_fu_3202;
reg   [15:0] tmp_V_450_fu_3206;
reg   [15:0] tmp_V_451_fu_3210;
reg   [15:0] tmp_V_452_fu_3214;
reg   [15:0] tmp_V_453_fu_3218;
reg   [15:0] tmp_V_454_fu_3222;
reg   [15:0] tmp_V_455_fu_3226;
reg   [15:0] tmp_V_456_fu_3230;
reg   [15:0] tmp_V_457_fu_3234;
reg   [15:0] tmp_V_458_fu_3238;
reg   [15:0] tmp_V_459_fu_3242;
reg   [15:0] tmp_V_460_fu_3246;
reg   [15:0] tmp_V_461_fu_3250;
reg   [15:0] tmp_V_462_fu_3254;
reg   [15:0] tmp_V_463_fu_3258;
reg   [15:0] tmp_V_464_fu_3262;
reg   [15:0] tmp_V_465_fu_3266;
reg   [15:0] tmp_V_466_fu_3270;
reg   [15:0] tmp_V_467_fu_3274;
reg   [15:0] tmp_V_468_fu_3278;
reg   [15:0] tmp_V_469_fu_3282;
reg   [15:0] tmp_V_470_fu_3286;
reg   [15:0] tmp_V_471_fu_3290;
reg   [15:0] tmp_V_472_fu_3294;
reg   [15:0] tmp_V_473_fu_3298;
reg   [15:0] tmp_V_474_fu_3302;
reg   [15:0] tmp_V_475_fu_3306;
reg   [15:0] tmp_V_476_fu_3310;
reg   [15:0] tmp_V_477_fu_3314;
reg   [15:0] tmp_V_478_fu_3318;
reg   [15:0] tmp_V_479_fu_3322;
reg   [15:0] tmp_V_480_fu_3326;
reg   [15:0] tmp_V_481_fu_3330;
reg   [15:0] tmp_V_482_fu_3334;
reg   [15:0] tmp_V_483_fu_3338;
reg   [15:0] tmp_V_484_fu_3342;
reg   [15:0] tmp_V_485_fu_3346;
reg   [15:0] tmp_V_486_fu_3350;
reg   [15:0] tmp_V_487_fu_3354;
reg   [15:0] tmp_V_488_fu_3358;
reg   [15:0] tmp_V_489_fu_3362;
reg   [15:0] tmp_V_490_fu_3366;
reg   [15:0] tmp_V_491_fu_3370;
reg   [15:0] tmp_V_492_fu_3374;
reg   [15:0] tmp_V_493_fu_3378;
reg   [15:0] tmp_V_494_fu_3382;
reg   [15:0] tmp_V_495_fu_3386;
reg   [15:0] tmp_V_496_fu_3390;
reg   [15:0] tmp_V_497_fu_3394;
reg   [15:0] tmp_V_498_fu_3398;
reg   [15:0] tmp_V_499_fu_3402;
reg   [15:0] tmp_V_500_fu_3406;
reg   [15:0] tmp_V_501_fu_3410;
reg   [15:0] tmp_V_502_fu_3414;
reg   [15:0] tmp_V_503_fu_3418;
reg   [15:0] tmp_V_504_fu_3422;
reg   [15:0] tmp_V_505_fu_3426;
reg   [15:0] tmp_V_506_fu_3430;
reg   [15:0] tmp_V_507_fu_3434;
reg   [15:0] tmp_V_508_fu_3438;
reg   [15:0] tmp_V_509_fu_3442;
reg   [15:0] tmp_V_510_fu_3446;
reg   [15:0] tmp_V_511_fu_3450;
reg   [15:0] tmp_V_512_fu_3454;
reg   [15:0] tmp_V_513_fu_3458;
reg   [15:0] tmp_V_514_fu_3462;
reg   [15:0] tmp_V_515_fu_3466;
reg   [15:0] tmp_V_516_fu_3470;
reg   [15:0] tmp_V_517_fu_3474;
reg   [15:0] tmp_V_518_fu_3478;
reg   [15:0] tmp_V_519_fu_3482;
reg   [15:0] tmp_V_520_fu_3486;
reg   [15:0] tmp_V_521_fu_3490;
reg   [15:0] tmp_V_522_fu_3494;
reg   [15:0] tmp_V_523_fu_3498;
reg   [15:0] tmp_V_524_fu_3502;
reg   [15:0] tmp_V_525_fu_3506;
reg   [15:0] tmp_V_526_fu_3510;
reg   [15:0] tmp_V_527_fu_3514;
reg   [15:0] tmp_V_528_fu_3518;
reg   [15:0] tmp_V_529_fu_3522;
reg   [15:0] tmp_V_530_fu_3526;
reg   [15:0] tmp_V_531_fu_3530;
reg   [15:0] tmp_V_532_fu_3534;
reg   [15:0] tmp_V_533_fu_3538;
reg   [15:0] tmp_V_534_fu_3542;
reg   [15:0] tmp_V_535_fu_3546;
reg   [15:0] tmp_V_536_fu_3550;
reg   [15:0] tmp_V_537_fu_3554;
reg   [15:0] tmp_V_538_fu_3558;
reg   [15:0] tmp_V_539_fu_3562;
reg   [15:0] tmp_V_540_fu_3566;
reg   [15:0] tmp_V_541_fu_3570;
reg   [15:0] tmp_V_542_fu_3574;
reg   [15:0] tmp_V_543_fu_3578;
reg   [15:0] tmp_V_544_fu_3582;
reg   [15:0] tmp_V_545_fu_3586;
reg   [15:0] tmp_V_546_fu_3590;
reg   [15:0] tmp_V_547_fu_3594;
reg   [15:0] tmp_V_548_fu_3598;
reg   [15:0] tmp_V_549_fu_3602;
reg   [15:0] tmp_V_550_fu_3606;
reg   [15:0] tmp_V_551_fu_3610;
reg   [15:0] tmp_V_552_fu_3614;
reg   [15:0] tmp_V_553_fu_3618;
reg   [15:0] tmp_V_554_fu_3622;
reg   [15:0] tmp_V_555_fu_3626;
reg   [15:0] tmp_V_556_fu_3630;
reg   [15:0] tmp_V_557_fu_3634;
reg   [15:0] tmp_V_558_fu_3638;
reg   [15:0] tmp_V_559_fu_3642;
reg   [15:0] tmp_V_560_fu_3646;
reg   [15:0] tmp_V_561_fu_3650;
reg   [15:0] tmp_V_562_fu_3654;
reg   [15:0] tmp_V_563_fu_3658;
reg   [15:0] tmp_V_564_fu_3662;
reg   [15:0] tmp_V_565_fu_3666;
reg   [15:0] tmp_V_566_fu_3670;
reg   [15:0] tmp_V_567_fu_3674;
reg   [15:0] tmp_V_568_fu_3678;
reg   [15:0] tmp_V_569_fu_3682;
reg   [15:0] tmp_V_570_fu_3686;
reg   [15:0] tmp_V_571_fu_3690;
reg   [15:0] tmp_V_572_fu_3694;
reg   [15:0] tmp_V_573_fu_3698;
reg   [15:0] tmp_V_574_fu_3702;
reg   [15:0] tmp_V_575_fu_3706;
reg   [15:0] tmp_V_576_fu_3710;
reg   [31:0] nf_assign_fu_3714;
wire   [31:0] select_ln301_fu_11988_p3;
reg   [31:0] ap_sig_allocacmp_nf_assign_load_1;
reg    ap_block_pp0_stage0_01001;
wire   [9:0] inElem_V_1_fu_7401_p577;
wire   [3:0] trunc_ln647_1_fu_11623_p1;
wire  signed [3:0] mul_ln1352_fu_11634_p0;
wire  signed [7:0] sext_ln215_1_fu_11630_p1;
wire  signed [7:0] mul_ln1352_fu_11634_p2;
wire   [3:0] arg_V_read_assign_1_fu_11644_p4;
wire  signed [3:0] mul_ln1352_1_fu_11661_p0;
wire  signed [7:0] sext_ln215_3_fu_11657_p1;
wire   [3:0] arg_V_read_assign_2_fu_11667_p4;
wire  signed [3:0] mul_ln1352_2_fu_11684_p0;
wire  signed [7:0] sext_ln215_5_fu_11680_p1;
wire  signed [7:0] mul_ln1352_2_fu_11684_p2;
wire   [3:0] arg_V_read_assign_3_fu_11694_p4;
wire  signed [3:0] mul_ln1352_3_fu_11711_p0;
wire  signed [7:0] sext_ln215_7_fu_11707_p1;
wire  signed [7:0] mul_ln1352_3_fu_11711_p2;
wire  signed [8:0] sext_ln700_1_fu_11717_p1;
wire  signed [8:0] sext_ln170_fu_11640_p1;
wire  signed [8:0] sext_ln170_1_fu_11690_p1;
wire   [8:0] add_ln700_1_fu_11721_p2;
wire  signed [3:0] mul_ln1352_4_fu_11736_p0;
wire  signed [7:0] mul_ln1352_4_fu_11736_p2;
wire  signed [3:0] mul_ln1352_5_fu_11749_p0;
wire  signed [3:0] mul_ln1352_6_fu_11758_p0;
wire  signed [7:0] mul_ln1352_6_fu_11758_p2;
wire  signed [3:0] mul_ln1352_7_fu_11771_p0;
wire  signed [7:0] mul_ln1352_7_fu_11771_p2;
wire  signed [8:0] sext_ln700_4_fu_11777_p1;
wire  signed [8:0] sext_ln170_2_fu_11742_p1;
wire  signed [8:0] sext_ln170_3_fu_11764_p1;
wire   [8:0] add_ln700_5_fu_11781_p2;
wire  signed [3:0] mul_ln1352_8_fu_11796_p0;
wire  signed [7:0] mul_ln1352_8_fu_11796_p2;
wire  signed [3:0] mul_ln1352_9_fu_11809_p0;
wire  signed [3:0] mul_ln1352_10_fu_11818_p0;
wire  signed [7:0] mul_ln1352_10_fu_11818_p2;
wire  signed [3:0] mul_ln1352_11_fu_11831_p0;
wire  signed [7:0] mul_ln1352_11_fu_11831_p2;
wire  signed [8:0] sext_ln700_7_fu_11837_p1;
wire  signed [8:0] sext_ln170_4_fu_11802_p1;
wire  signed [8:0] sext_ln170_5_fu_11824_p1;
wire   [8:0] add_ln700_9_fu_11841_p2;
wire  signed [3:0] mul_ln1352_12_fu_11856_p0;
wire  signed [7:0] mul_ln1352_12_fu_11856_p2;
wire  signed [3:0] mul_ln1352_13_fu_11869_p0;
wire  signed [3:0] mul_ln1352_14_fu_11878_p0;
wire  signed [7:0] mul_ln1352_14_fu_11878_p2;
wire  signed [3:0] mul_ln1352_15_fu_11891_p0;
wire  signed [7:0] mul_ln1352_15_fu_11891_p2;
wire  signed [8:0] sext_ln700_10_fu_11897_p1;
wire  signed [8:0] sext_ln170_6_fu_11862_p1;
wire  signed [8:0] sext_ln170_7_fu_11884_p1;
wire   [8:0] add_ln700_13_fu_11901_p2;
wire   [31:0] nf_fu_11976_p2;
wire   [0:0] icmp_ln301_fu_11982_p2;
wire  signed [17:0] sext_ln700_fu_12041_p1;
wire   [17:0] select_ln271_3_fu_12034_p3;
wire   [17:0] add_ln700_fu_12044_p2;
wire  signed [17:0] sext_ln700_2_fu_12050_p1;
wire  signed [17:0] sext_ln700_3_fu_12059_p1;
wire   [17:0] select_ln271_2_fu_12027_p3;
wire   [17:0] add_ln700_4_fu_12062_p2;
wire  signed [17:0] sext_ln700_5_fu_12068_p1;
wire  signed [17:0] sext_ln700_6_fu_12077_p1;
wire   [17:0] select_ln271_1_fu_12020_p3;
wire   [17:0] add_ln700_8_fu_12080_p2;
wire  signed [17:0] sext_ln700_8_fu_12086_p1;
wire  signed [17:0] sext_ln700_9_fu_12095_p1;
wire   [17:0] select_ln271_fu_12013_p3;
wire   [17:0] add_ln700_12_fu_12098_p2;
wire  signed [17:0] sext_ln700_11_fu_12104_p1;
wire  signed [17:0] sext_ln142_fu_12133_p1;
wire  signed [17:0] sext_ln142_1_fu_12143_p1;
wire  signed [17:0] sext_ln142_2_fu_12153_p1;
wire  signed [17:0] sext_ln142_3_fu_12163_p1;
wire  signed [17:0] sext_ln142_4_fu_12173_p1;
wire  signed [17:0] sext_ln142_5_fu_12183_p1;
wire  signed [17:0] sext_ln142_6_fu_12193_p1;
wire  signed [17:0] sext_ln142_7_fu_12203_p1;
wire  signed [17:0] sext_ln142_8_fu_12213_p1;
wire  signed [17:0] sext_ln142_9_fu_12223_p1;
wire  signed [17:0] sext_ln142_10_fu_12233_p1;
wire  signed [17:0] sext_ln142_11_fu_12243_p1;
wire  signed [17:0] sext_ln142_12_fu_12253_p1;
wire  signed [17:0] sext_ln142_13_fu_12263_p1;
wire  signed [17:0] sext_ln142_14_fu_12357_p1;
wire  signed [17:0] sext_ln142_15_fu_12367_p1;
wire  signed [17:0] sext_ln142_16_fu_12377_p1;
wire  signed [17:0] sext_ln142_17_fu_12387_p1;
wire  signed [17:0] sext_ln142_18_fu_12397_p1;
wire  signed [17:0] sext_ln142_19_fu_12407_p1;
wire  signed [17:0] sext_ln142_20_fu_12417_p1;
wire  signed [17:0] sext_ln142_21_fu_12427_p1;
wire  signed [17:0] sext_ln142_22_fu_12437_p1;
wire  signed [17:0] sext_ln142_23_fu_12447_p1;
wire  signed [17:0] sext_ln142_24_fu_12457_p1;
wire  signed [17:0] sext_ln142_25_fu_12467_p1;
wire  signed [17:0] sext_ln142_26_fu_12477_p1;
wire  signed [17:0] sext_ln142_27_fu_12487_p1;
wire  signed [17:0] sext_ln142_28_fu_12503_p1;
wire  signed [17:0] sext_ln142_29_fu_12513_p1;
wire  signed [17:0] sext_ln142_30_fu_12523_p1;
wire  signed [17:0] sext_ln142_31_fu_12533_p1;
wire  signed [17:0] sext_ln142_32_fu_12543_p1;
wire  signed [17:0] sext_ln142_33_fu_12553_p1;
wire  signed [17:0] sext_ln142_34_fu_12563_p1;
wire  signed [17:0] sext_ln142_35_fu_12573_p1;
wire  signed [17:0] sext_ln142_36_fu_12583_p1;
wire  signed [17:0] sext_ln142_37_fu_12593_p1;
wire  signed [17:0] sext_ln142_38_fu_12603_p1;
wire   [0:0] xor_ln899_fu_12625_p2;
wire   [0:0] xor_ln899_1_fu_12634_p2;
wire   [0:0] xor_ln899_2_fu_12643_p2;
wire   [0:0] xor_ln899_3_fu_12652_p2;
wire   [0:0] xor_ln899_4_fu_12661_p2;
wire   [0:0] xor_ln899_5_fu_12670_p2;
wire   [0:0] xor_ln899_6_fu_12679_p2;
wire   [0:0] xor_ln899_7_fu_12688_p2;
wire   [0:0] xor_ln899_8_fu_12697_p2;
wire   [0:0] xor_ln899_9_fu_12706_p2;
wire   [0:0] xor_ln899_10_fu_12715_p2;
wire   [0:0] xor_ln899_11_fu_12724_p2;
wire   [0:0] xor_ln899_12_fu_12733_p2;
wire   [0:0] xor_ln899_13_fu_12742_p2;
wire   [1:0] zext_ln142_2_fu_12639_p1;
wire   [1:0] zext_ln142_3_fu_12648_p1;
wire   [1:0] add_ln700_16_fu_12751_p2;
wire   [1:0] zext_ln142_1_fu_12630_p1;
wire   [1:0] add_ln700_17_fu_12757_p2;
wire   [1:0] zext_ln142_4_fu_12657_p1;
wire   [1:0] zext_ln142_5_fu_12666_p1;
wire   [1:0] add_ln700_18_fu_12767_p2;
wire   [1:0] zext_ln142_6_fu_12675_p1;
wire   [1:0] zext_ln142_7_fu_12684_p1;
wire   [1:0] add_ln700_19_fu_12777_p2;
wire   [2:0] zext_ln700_3_fu_12783_p1;
wire   [2:0] zext_ln700_2_fu_12773_p1;
wire   [2:0] add_ln700_20_fu_12787_p2;
wire   [2:0] zext_ln700_1_fu_12763_p1;
wire   [2:0] add_ln700_21_fu_12793_p2;
wire   [1:0] zext_ln142_9_fu_12702_p1;
wire   [1:0] zext_ln142_10_fu_12711_p1;
wire   [1:0] add_ln700_22_fu_12803_p2;
wire   [1:0] zext_ln142_8_fu_12693_p1;
wire   [1:0] add_ln700_23_fu_12809_p2;
wire   [1:0] zext_ln142_11_fu_12720_p1;
wire   [1:0] zext_ln142_12_fu_12729_p1;
wire   [1:0] add_ln700_24_fu_12819_p2;
wire   [1:0] zext_ln142_13_fu_12738_p1;
wire   [1:0] zext_ln700_fu_12747_p1;
wire   [1:0] add_ln700_25_fu_12829_p2;
wire   [2:0] zext_ln700_7_fu_12835_p1;
wire   [2:0] zext_ln700_6_fu_12825_p1;
wire   [2:0] add_ln700_26_fu_12839_p2;
wire   [2:0] zext_ln700_5_fu_12815_p1;
wire   [2:0] add_ln700_27_fu_12845_p2;
wire   [3:0] zext_ln700_8_fu_12851_p1;
wire   [3:0] zext_ln700_4_fu_12799_p1;
wire   [0:0] xor_ln899_14_fu_12861_p2;
wire   [0:0] xor_ln899_15_fu_12870_p2;
wire   [0:0] xor_ln899_16_fu_12879_p2;
wire   [0:0] xor_ln899_17_fu_12888_p2;
wire   [0:0] xor_ln899_18_fu_12897_p2;
wire   [0:0] xor_ln899_19_fu_12906_p2;
wire   [0:0] xor_ln899_20_fu_12915_p2;
wire   [0:0] xor_ln899_21_fu_12924_p2;
wire   [0:0] xor_ln899_22_fu_12933_p2;
wire   [0:0] xor_ln899_23_fu_12942_p2;
wire   [0:0] xor_ln899_24_fu_12951_p2;
wire   [0:0] xor_ln899_25_fu_12960_p2;
wire   [0:0] xor_ln899_26_fu_12969_p2;
wire   [0:0] xor_ln899_27_fu_12978_p2;
wire   [1:0] zext_ln142_15_fu_12875_p1;
wire   [1:0] zext_ln142_16_fu_12884_p1;
wire   [1:0] add_ln700_29_fu_12987_p2;
wire   [1:0] zext_ln142_14_fu_12866_p1;
wire   [1:0] add_ln700_30_fu_12993_p2;
wire   [1:0] zext_ln142_17_fu_12893_p1;
wire   [1:0] zext_ln142_18_fu_12902_p1;
wire   [1:0] add_ln700_31_fu_13003_p2;
wire   [1:0] zext_ln142_19_fu_12911_p1;
wire   [1:0] zext_ln142_20_fu_12920_p1;
wire   [1:0] add_ln700_32_fu_13013_p2;
wire   [2:0] zext_ln700_12_fu_13019_p1;
wire   [2:0] zext_ln700_11_fu_13009_p1;
wire   [2:0] add_ln700_33_fu_13023_p2;
wire   [2:0] zext_ln700_10_fu_12999_p1;
wire   [2:0] add_ln700_34_fu_13029_p2;
wire   [1:0] zext_ln142_22_fu_12938_p1;
wire   [1:0] zext_ln142_23_fu_12947_p1;
wire   [1:0] add_ln700_35_fu_13039_p2;
wire   [1:0] zext_ln142_21_fu_12929_p1;
wire   [1:0] add_ln700_36_fu_13045_p2;
wire   [1:0] zext_ln142_24_fu_12956_p1;
wire   [1:0] zext_ln142_25_fu_12965_p1;
wire   [1:0] add_ln700_37_fu_13055_p2;
wire   [1:0] zext_ln142_26_fu_12974_p1;
wire   [1:0] zext_ln700_9_fu_12983_p1;
wire   [1:0] add_ln700_38_fu_13065_p2;
wire   [2:0] zext_ln700_16_fu_13071_p1;
wire   [2:0] zext_ln700_15_fu_13061_p1;
wire   [2:0] add_ln700_39_fu_13075_p2;
wire   [2:0] zext_ln700_14_fu_13051_p1;
wire   [2:0] add_ln700_40_fu_13081_p2;
wire   [3:0] zext_ln700_17_fu_13087_p1;
wire   [3:0] zext_ln700_13_fu_13035_p1;
wire   [0:0] xor_ln899_28_fu_13097_p2;
wire   [0:0] xor_ln899_29_fu_13106_p2;
wire   [0:0] xor_ln899_30_fu_13115_p2;
wire   [0:0] xor_ln899_31_fu_13124_p2;
wire   [0:0] xor_ln899_32_fu_13133_p2;
wire   [0:0] xor_ln899_33_fu_13142_p2;
wire   [0:0] xor_ln899_34_fu_13151_p2;
wire   [0:0] xor_ln899_35_fu_13160_p2;
wire   [0:0] xor_ln899_36_fu_13169_p2;
wire   [0:0] xor_ln899_37_fu_13178_p2;
wire   [0:0] xor_ln899_38_fu_13187_p2;
wire   [0:0] xor_ln899_39_fu_13196_p2;
wire   [0:0] xor_ln899_40_fu_13205_p2;
wire   [0:0] xor_ln899_41_fu_13214_p2;
wire   [1:0] zext_ln142_28_fu_13111_p1;
wire   [1:0] zext_ln142_29_fu_13120_p1;
wire   [1:0] add_ln700_42_fu_13223_p2;
wire   [1:0] zext_ln142_27_fu_13102_p1;
wire   [1:0] add_ln700_43_fu_13229_p2;
wire   [1:0] zext_ln142_30_fu_13129_p1;
wire   [1:0] zext_ln142_31_fu_13138_p1;
wire   [1:0] add_ln700_44_fu_13239_p2;
wire   [1:0] zext_ln142_32_fu_13147_p1;
wire   [1:0] zext_ln142_33_fu_13156_p1;
wire   [1:0] add_ln700_45_fu_13249_p2;
wire   [2:0] zext_ln700_21_fu_13255_p1;
wire   [2:0] zext_ln700_20_fu_13245_p1;
wire   [2:0] add_ln700_46_fu_13259_p2;
wire   [2:0] zext_ln700_19_fu_13235_p1;
wire   [2:0] add_ln700_47_fu_13265_p2;
wire   [1:0] zext_ln142_35_fu_13174_p1;
wire   [1:0] zext_ln142_36_fu_13183_p1;
wire   [1:0] add_ln700_48_fu_13275_p2;
wire   [1:0] zext_ln142_34_fu_13165_p1;
wire   [1:0] add_ln700_49_fu_13281_p2;
wire   [1:0] zext_ln142_37_fu_13192_p1;
wire   [1:0] zext_ln142_38_fu_13201_p1;
wire   [1:0] add_ln700_50_fu_13291_p2;
wire   [1:0] zext_ln142_39_fu_13210_p1;
wire   [1:0] zext_ln700_18_fu_13219_p1;
wire   [1:0] add_ln700_51_fu_13301_p2;
wire   [2:0] zext_ln700_25_fu_13307_p1;
wire   [2:0] zext_ln700_24_fu_13297_p1;
wire   [2:0] add_ln700_52_fu_13311_p2;
wire   [2:0] zext_ln700_23_fu_13287_p1;
wire   [2:0] add_ln700_53_fu_13317_p2;
wire   [3:0] zext_ln700_26_fu_13323_p1;
wire   [3:0] zext_ln700_22_fu_13271_p1;
wire   [0:0] xor_ln899_42_fu_13333_p2;
wire   [0:0] xor_ln899_43_fu_13342_p2;
wire   [0:0] xor_ln899_44_fu_13351_p2;
wire   [0:0] xor_ln899_45_fu_13360_p2;
wire   [0:0] xor_ln899_46_fu_13369_p2;
wire   [0:0] xor_ln899_47_fu_13378_p2;
wire   [0:0] xor_ln899_48_fu_13387_p2;
wire   [0:0] xor_ln899_49_fu_13396_p2;
wire   [0:0] xor_ln899_50_fu_13405_p2;
wire   [0:0] xor_ln899_51_fu_13414_p2;
wire   [0:0] xor_ln899_52_fu_13423_p2;
wire   [0:0] xor_ln899_53_fu_13432_p2;
wire   [0:0] xor_ln899_54_fu_13441_p2;
wire   [0:0] xor_ln899_55_fu_13450_p2;
wire   [1:0] zext_ln142_41_fu_13347_p1;
wire   [1:0] zext_ln142_42_fu_13356_p1;
wire   [1:0] add_ln700_55_fu_13459_p2;
wire   [1:0] zext_ln142_40_fu_13338_p1;
wire   [1:0] add_ln700_56_fu_13465_p2;
wire   [1:0] zext_ln142_43_fu_13365_p1;
wire   [1:0] zext_ln142_44_fu_13374_p1;
wire   [1:0] add_ln700_57_fu_13475_p2;
wire   [1:0] zext_ln142_45_fu_13383_p1;
wire   [1:0] zext_ln142_46_fu_13392_p1;
wire   [1:0] add_ln700_58_fu_13485_p2;
wire   [2:0] zext_ln700_30_fu_13491_p1;
wire   [2:0] zext_ln700_29_fu_13481_p1;
wire   [2:0] add_ln700_59_fu_13495_p2;
wire   [2:0] zext_ln700_28_fu_13471_p1;
wire   [2:0] add_ln700_60_fu_13501_p2;
wire   [1:0] zext_ln142_48_fu_13410_p1;
wire   [1:0] zext_ln142_49_fu_13419_p1;
wire   [1:0] add_ln700_61_fu_13511_p2;
wire   [1:0] zext_ln142_47_fu_13401_p1;
wire   [1:0] add_ln700_62_fu_13517_p2;
wire   [1:0] zext_ln142_50_fu_13428_p1;
wire   [1:0] zext_ln142_51_fu_13437_p1;
wire   [1:0] add_ln700_63_fu_13527_p2;
wire   [1:0] zext_ln142_52_fu_13446_p1;
wire   [1:0] zext_ln700_27_fu_13455_p1;
wire   [1:0] add_ln700_64_fu_13537_p2;
wire   [2:0] zext_ln700_34_fu_13543_p1;
wire   [2:0] zext_ln700_33_fu_13533_p1;
wire   [2:0] add_ln700_65_fu_13547_p2;
wire   [2:0] zext_ln700_32_fu_13523_p1;
wire   [2:0] add_ln700_66_fu_13553_p2;
wire   [3:0] zext_ln700_35_fu_13559_p1;
wire   [3:0] zext_ln700_31_fu_13507_p1;
wire   [3:0] add_ln700_67_fu_13563_p2;
wire   [3:0] add_ln700_54_fu_13327_p2;
wire   [3:0] add_ln700_41_fu_13091_p2;
wire   [3:0] add_ln700_28_fu_12855_p2;
wire    ap_CS_fsm_state6;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

StreamingFCLayer_Batch_1_Matrix_Vector_Actbkb #(
    .DataWidth( 16 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_55_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_55_address0),
    .ce0(threshs_m_thresholds_55_ce0),
    .q0(threshs_m_thresholds_55_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actcud #(
    .DataWidth( 16 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_54_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_54_address0),
    .ce0(threshs_m_thresholds_54_ce0),
    .q0(threshs_m_thresholds_54_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActdEe #(
    .DataWidth( 16 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_49_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_49_address0),
    .ce0(threshs_m_thresholds_49_ce0),
    .q0(threshs_m_thresholds_49_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActeOg #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_48_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_48_address0),
    .ce0(threshs_m_thresholds_48_ce0),
    .q0(threshs_m_thresholds_48_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActfYi #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_47_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_47_address0),
    .ce0(threshs_m_thresholds_47_ce0),
    .q0(threshs_m_thresholds_47_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actg8j #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_46_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_46_address0),
    .ce0(threshs_m_thresholds_46_ce0),
    .q0(threshs_m_thresholds_46_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Acthbi #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_45_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_45_address0),
    .ce0(threshs_m_thresholds_45_ce0),
    .q0(threshs_m_thresholds_45_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actibs #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_44_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_44_address0),
    .ce0(threshs_m_thresholds_44_ce0),
    .q0(threshs_m_thresholds_44_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActjbC #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_43_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_43_address0),
    .ce0(threshs_m_thresholds_43_ce0),
    .q0(threshs_m_thresholds_43_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActkbM #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_42_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_42_address0),
    .ce0(threshs_m_thresholds_42_ce0),
    .q0(threshs_m_thresholds_42_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActlbW #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_53_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_53_address0),
    .ce0(threshs_m_thresholds_53_ce0),
    .q0(threshs_m_thresholds_53_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actmb6 #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_52_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_52_address0),
    .ce0(threshs_m_thresholds_52_ce0),
    .q0(threshs_m_thresholds_52_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actncg #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_51_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_51_address0),
    .ce0(threshs_m_thresholds_51_ce0),
    .q0(threshs_m_thresholds_51_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actocq #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_50_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_50_address0),
    .ce0(threshs_m_thresholds_50_ce0),
    .q0(threshs_m_thresholds_50_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActpcA #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_41_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_41_address0),
    .ce0(threshs_m_thresholds_41_ce0),
    .q0(threshs_m_thresholds_41_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActqcK #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_40_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_40_address0),
    .ce0(threshs_m_thresholds_40_ce0),
    .q0(threshs_m_thresholds_40_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActrcU #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_35_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_35_address0),
    .ce0(threshs_m_thresholds_35_ce0),
    .q0(threshs_m_thresholds_35_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actsc4 #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_34_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_34_address0),
    .ce0(threshs_m_thresholds_34_ce0),
    .q0(threshs_m_thresholds_34_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Acttde #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_33_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_33_address0),
    .ce0(threshs_m_thresholds_33_ce0),
    .q0(threshs_m_thresholds_33_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actudo #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_32_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_32_address0),
    .ce0(threshs_m_thresholds_32_ce0),
    .q0(threshs_m_thresholds_32_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actvdy #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_31_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_31_address0),
    .ce0(threshs_m_thresholds_31_ce0),
    .q0(threshs_m_thresholds_31_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActwdI #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_30_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_30_address0),
    .ce0(threshs_m_thresholds_30_ce0),
    .q0(threshs_m_thresholds_30_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActxdS #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_29_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_29_address0),
    .ce0(threshs_m_thresholds_29_ce0),
    .q0(threshs_m_thresholds_29_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actyd2 #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_28_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_28_address0),
    .ce0(threshs_m_thresholds_28_ce0),
    .q0(threshs_m_thresholds_28_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Actzec #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_39_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_39_address0),
    .ce0(threshs_m_thresholds_39_ce0),
    .q0(threshs_m_thresholds_39_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActAem #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_38_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_38_address0),
    .ce0(threshs_m_thresholds_38_ce0),
    .q0(threshs_m_thresholds_38_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActBew #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_37_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_37_address0),
    .ce0(threshs_m_thresholds_37_ce0),
    .q0(threshs_m_thresholds_37_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActCeG #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_36_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_36_address0),
    .ce0(threshs_m_thresholds_36_ce0),
    .q0(threshs_m_thresholds_36_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActDeQ #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_27_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_27_address0),
    .ce0(threshs_m_thresholds_27_ce0),
    .q0(threshs_m_thresholds_27_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActEe0 #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_26_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_26_address0),
    .ce0(threshs_m_thresholds_26_ce0),
    .q0(threshs_m_thresholds_26_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActFfa #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_21_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_21_address0),
    .ce0(threshs_m_thresholds_21_ce0),
    .q0(threshs_m_thresholds_21_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActGfk #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_20_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_20_address0),
    .ce0(threshs_m_thresholds_20_ce0),
    .q0(threshs_m_thresholds_20_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActHfu #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_19_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_19_address0),
    .ce0(threshs_m_thresholds_19_ce0),
    .q0(threshs_m_thresholds_19_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActIfE #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_18_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_18_address0),
    .ce0(threshs_m_thresholds_18_ce0),
    .q0(threshs_m_thresholds_18_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActJfO #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_17_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_17_address0),
    .ce0(threshs_m_thresholds_17_ce0),
    .q0(threshs_m_thresholds_17_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActKfY #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_16_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_16_address0),
    .ce0(threshs_m_thresholds_16_ce0),
    .q0(threshs_m_thresholds_16_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActLf8 #(
    .DataWidth( 16 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_15_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_15_address0),
    .ce0(threshs_m_thresholds_15_ce0),
    .q0(threshs_m_thresholds_15_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActMgi #(
    .DataWidth( 16 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_14_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_14_address0),
    .ce0(threshs_m_thresholds_14_ce0),
    .q0(threshs_m_thresholds_14_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActNgs #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_25_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_25_address0),
    .ce0(threshs_m_thresholds_25_ce0),
    .q0(threshs_m_thresholds_25_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActOgC #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_24_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_24_address0),
    .ce0(threshs_m_thresholds_24_ce0),
    .q0(threshs_m_thresholds_24_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActPgM #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_23_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_23_address0),
    .ce0(threshs_m_thresholds_23_ce0),
    .q0(threshs_m_thresholds_23_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActQgW #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_22_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_22_address0),
    .ce0(threshs_m_thresholds_22_ce0),
    .q0(threshs_m_thresholds_22_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActRg6 #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_13_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_13_address0),
    .ce0(threshs_m_thresholds_13_ce0),
    .q0(threshs_m_thresholds_13_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActShg #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_12_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_12_address0),
    .ce0(threshs_m_thresholds_12_ce0),
    .q0(threshs_m_thresholds_12_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActThq #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_7_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_7_address0),
    .ce0(threshs_m_thresholds_7_ce0),
    .q0(threshs_m_thresholds_7_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActUhA #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_6_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_6_address0),
    .ce0(threshs_m_thresholds_6_ce0),
    .q0(threshs_m_thresholds_6_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActVhK #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_5_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_5_address0),
    .ce0(threshs_m_thresholds_5_ce0),
    .q0(threshs_m_thresholds_5_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActWhU #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_4_address0),
    .ce0(threshs_m_thresholds_4_ce0),
    .q0(threshs_m_thresholds_4_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActXh4 #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_3_address0),
    .ce0(threshs_m_thresholds_3_ce0),
    .q0(threshs_m_thresholds_3_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActYie #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_2_address0),
    .ce0(threshs_m_thresholds_2_ce0),
    .q0(threshs_m_thresholds_2_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_ActZio #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_1_address0),
    .ce0(threshs_m_thresholds_1_ce0),
    .q0(threshs_m_thresholds_1_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Act0iy #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_address0),
    .ce0(threshs_m_thresholds_ce0),
    .q0(threshs_m_thresholds_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Act1iI #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_11_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_11_address0),
    .ce0(threshs_m_thresholds_11_ce0),
    .q0(threshs_m_thresholds_11_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Act2iS #(
    .DataWidth( 17 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_10_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_10_address0),
    .ce0(threshs_m_thresholds_10_ce0),
    .q0(threshs_m_thresholds_10_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Act3i2 #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_9_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_9_address0),
    .ce0(threshs_m_thresholds_9_ce0),
    .q0(threshs_m_thresholds_9_q0)
);

StreamingFCLayer_Batch_1_Matrix_Vector_Act4jc #(
    .DataWidth( 18 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
threshs_m_thresholds_8_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_8_address0),
    .ce0(threshs_m_thresholds_8_ce0),
    .q0(threshs_m_thresholds_8_q0)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_5jm #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .din2_WIDTH( 16 ),
    .din3_WIDTH( 16 ),
    .din4_WIDTH( 16 ),
    .din5_WIDTH( 16 ),
    .din6_WIDTH( 16 ),
    .din7_WIDTH( 16 ),
    .din8_WIDTH( 16 ),
    .din9_WIDTH( 16 ),
    .din10_WIDTH( 16 ),
    .din11_WIDTH( 16 ),
    .din12_WIDTH( 16 ),
    .din13_WIDTH( 16 ),
    .din14_WIDTH( 16 ),
    .din15_WIDTH( 16 ),
    .din16_WIDTH( 16 ),
    .din17_WIDTH( 16 ),
    .din18_WIDTH( 16 ),
    .din19_WIDTH( 16 ),
    .din20_WIDTH( 16 ),
    .din21_WIDTH( 16 ),
    .din22_WIDTH( 16 ),
    .din23_WIDTH( 16 ),
    .din24_WIDTH( 16 ),
    .din25_WIDTH( 16 ),
    .din26_WIDTH( 16 ),
    .din27_WIDTH( 16 ),
    .din28_WIDTH( 16 ),
    .din29_WIDTH( 16 ),
    .din30_WIDTH( 16 ),
    .din31_WIDTH( 16 ),
    .din32_WIDTH( 16 ),
    .din33_WIDTH( 16 ),
    .din34_WIDTH( 16 ),
    .din35_WIDTH( 16 ),
    .din36_WIDTH( 16 ),
    .din37_WIDTH( 16 ),
    .din38_WIDTH( 16 ),
    .din39_WIDTH( 16 ),
    .din40_WIDTH( 16 ),
    .din41_WIDTH( 16 ),
    .din42_WIDTH( 16 ),
    .din43_WIDTH( 16 ),
    .din44_WIDTH( 16 ),
    .din45_WIDTH( 16 ),
    .din46_WIDTH( 16 ),
    .din47_WIDTH( 16 ),
    .din48_WIDTH( 16 ),
    .din49_WIDTH( 16 ),
    .din50_WIDTH( 16 ),
    .din51_WIDTH( 16 ),
    .din52_WIDTH( 16 ),
    .din53_WIDTH( 16 ),
    .din54_WIDTH( 16 ),
    .din55_WIDTH( 16 ),
    .din56_WIDTH( 16 ),
    .din57_WIDTH( 16 ),
    .din58_WIDTH( 16 ),
    .din59_WIDTH( 16 ),
    .din60_WIDTH( 16 ),
    .din61_WIDTH( 16 ),
    .din62_WIDTH( 16 ),
    .din63_WIDTH( 16 ),
    .din64_WIDTH( 16 ),
    .din65_WIDTH( 16 ),
    .din66_WIDTH( 16 ),
    .din67_WIDTH( 16 ),
    .din68_WIDTH( 16 ),
    .din69_WIDTH( 16 ),
    .din70_WIDTH( 16 ),
    .din71_WIDTH( 16 ),
    .din72_WIDTH( 16 ),
    .din73_WIDTH( 16 ),
    .din74_WIDTH( 16 ),
    .din75_WIDTH( 16 ),
    .din76_WIDTH( 16 ),
    .din77_WIDTH( 16 ),
    .din78_WIDTH( 16 ),
    .din79_WIDTH( 16 ),
    .din80_WIDTH( 16 ),
    .din81_WIDTH( 16 ),
    .din82_WIDTH( 16 ),
    .din83_WIDTH( 16 ),
    .din84_WIDTH( 16 ),
    .din85_WIDTH( 16 ),
    .din86_WIDTH( 16 ),
    .din87_WIDTH( 16 ),
    .din88_WIDTH( 16 ),
    .din89_WIDTH( 16 ),
    .din90_WIDTH( 16 ),
    .din91_WIDTH( 16 ),
    .din92_WIDTH( 16 ),
    .din93_WIDTH( 16 ),
    .din94_WIDTH( 16 ),
    .din95_WIDTH( 16 ),
    .din96_WIDTH( 16 ),
    .din97_WIDTH( 16 ),
    .din98_WIDTH( 16 ),
    .din99_WIDTH( 16 ),
    .din100_WIDTH( 16 ),
    .din101_WIDTH( 16 ),
    .din102_WIDTH( 16 ),
    .din103_WIDTH( 16 ),
    .din104_WIDTH( 16 ),
    .din105_WIDTH( 16 ),
    .din106_WIDTH( 16 ),
    .din107_WIDTH( 16 ),
    .din108_WIDTH( 16 ),
    .din109_WIDTH( 16 ),
    .din110_WIDTH( 16 ),
    .din111_WIDTH( 16 ),
    .din112_WIDTH( 16 ),
    .din113_WIDTH( 16 ),
    .din114_WIDTH( 16 ),
    .din115_WIDTH( 16 ),
    .din116_WIDTH( 16 ),
    .din117_WIDTH( 16 ),
    .din118_WIDTH( 16 ),
    .din119_WIDTH( 16 ),
    .din120_WIDTH( 16 ),
    .din121_WIDTH( 16 ),
    .din122_WIDTH( 16 ),
    .din123_WIDTH( 16 ),
    .din124_WIDTH( 16 ),
    .din125_WIDTH( 16 ),
    .din126_WIDTH( 16 ),
    .din127_WIDTH( 16 ),
    .din128_WIDTH( 16 ),
    .din129_WIDTH( 16 ),
    .din130_WIDTH( 16 ),
    .din131_WIDTH( 16 ),
    .din132_WIDTH( 16 ),
    .din133_WIDTH( 16 ),
    .din134_WIDTH( 16 ),
    .din135_WIDTH( 16 ),
    .din136_WIDTH( 16 ),
    .din137_WIDTH( 16 ),
    .din138_WIDTH( 16 ),
    .din139_WIDTH( 16 ),
    .din140_WIDTH( 16 ),
    .din141_WIDTH( 16 ),
    .din142_WIDTH( 16 ),
    .din143_WIDTH( 16 ),
    .din144_WIDTH( 16 ),
    .din145_WIDTH( 16 ),
    .din146_WIDTH( 16 ),
    .din147_WIDTH( 16 ),
    .din148_WIDTH( 16 ),
    .din149_WIDTH( 16 ),
    .din150_WIDTH( 16 ),
    .din151_WIDTH( 16 ),
    .din152_WIDTH( 16 ),
    .din153_WIDTH( 16 ),
    .din154_WIDTH( 16 ),
    .din155_WIDTH( 16 ),
    .din156_WIDTH( 16 ),
    .din157_WIDTH( 16 ),
    .din158_WIDTH( 16 ),
    .din159_WIDTH( 16 ),
    .din160_WIDTH( 16 ),
    .din161_WIDTH( 16 ),
    .din162_WIDTH( 16 ),
    .din163_WIDTH( 16 ),
    .din164_WIDTH( 16 ),
    .din165_WIDTH( 16 ),
    .din166_WIDTH( 16 ),
    .din167_WIDTH( 16 ),
    .din168_WIDTH( 16 ),
    .din169_WIDTH( 16 ),
    .din170_WIDTH( 16 ),
    .din171_WIDTH( 16 ),
    .din172_WIDTH( 16 ),
    .din173_WIDTH( 16 ),
    .din174_WIDTH( 16 ),
    .din175_WIDTH( 16 ),
    .din176_WIDTH( 16 ),
    .din177_WIDTH( 16 ),
    .din178_WIDTH( 16 ),
    .din179_WIDTH( 16 ),
    .din180_WIDTH( 16 ),
    .din181_WIDTH( 16 ),
    .din182_WIDTH( 16 ),
    .din183_WIDTH( 16 ),
    .din184_WIDTH( 16 ),
    .din185_WIDTH( 16 ),
    .din186_WIDTH( 16 ),
    .din187_WIDTH( 16 ),
    .din188_WIDTH( 16 ),
    .din189_WIDTH( 16 ),
    .din190_WIDTH( 16 ),
    .din191_WIDTH( 16 ),
    .din192_WIDTH( 16 ),
    .din193_WIDTH( 16 ),
    .din194_WIDTH( 16 ),
    .din195_WIDTH( 16 ),
    .din196_WIDTH( 16 ),
    .din197_WIDTH( 16 ),
    .din198_WIDTH( 16 ),
    .din199_WIDTH( 16 ),
    .din200_WIDTH( 16 ),
    .din201_WIDTH( 16 ),
    .din202_WIDTH( 16 ),
    .din203_WIDTH( 16 ),
    .din204_WIDTH( 16 ),
    .din205_WIDTH( 16 ),
    .din206_WIDTH( 16 ),
    .din207_WIDTH( 16 ),
    .din208_WIDTH( 16 ),
    .din209_WIDTH( 16 ),
    .din210_WIDTH( 16 ),
    .din211_WIDTH( 16 ),
    .din212_WIDTH( 16 ),
    .din213_WIDTH( 16 ),
    .din214_WIDTH( 16 ),
    .din215_WIDTH( 16 ),
    .din216_WIDTH( 16 ),
    .din217_WIDTH( 16 ),
    .din218_WIDTH( 16 ),
    .din219_WIDTH( 16 ),
    .din220_WIDTH( 16 ),
    .din221_WIDTH( 16 ),
    .din222_WIDTH( 16 ),
    .din223_WIDTH( 16 ),
    .din224_WIDTH( 16 ),
    .din225_WIDTH( 16 ),
    .din226_WIDTH( 16 ),
    .din227_WIDTH( 16 ),
    .din228_WIDTH( 16 ),
    .din229_WIDTH( 16 ),
    .din230_WIDTH( 16 ),
    .din231_WIDTH( 16 ),
    .din232_WIDTH( 16 ),
    .din233_WIDTH( 16 ),
    .din234_WIDTH( 16 ),
    .din235_WIDTH( 16 ),
    .din236_WIDTH( 16 ),
    .din237_WIDTH( 16 ),
    .din238_WIDTH( 16 ),
    .din239_WIDTH( 16 ),
    .din240_WIDTH( 16 ),
    .din241_WIDTH( 16 ),
    .din242_WIDTH( 16 ),
    .din243_WIDTH( 16 ),
    .din244_WIDTH( 16 ),
    .din245_WIDTH( 16 ),
    .din246_WIDTH( 16 ),
    .din247_WIDTH( 16 ),
    .din248_WIDTH( 16 ),
    .din249_WIDTH( 16 ),
    .din250_WIDTH( 16 ),
    .din251_WIDTH( 16 ),
    .din252_WIDTH( 16 ),
    .din253_WIDTH( 16 ),
    .din254_WIDTH( 16 ),
    .din255_WIDTH( 16 ),
    .din256_WIDTH( 16 ),
    .din257_WIDTH( 16 ),
    .din258_WIDTH( 16 ),
    .din259_WIDTH( 16 ),
    .din260_WIDTH( 16 ),
    .din261_WIDTH( 16 ),
    .din262_WIDTH( 16 ),
    .din263_WIDTH( 16 ),
    .din264_WIDTH( 16 ),
    .din265_WIDTH( 16 ),
    .din266_WIDTH( 16 ),
    .din267_WIDTH( 16 ),
    .din268_WIDTH( 16 ),
    .din269_WIDTH( 16 ),
    .din270_WIDTH( 16 ),
    .din271_WIDTH( 16 ),
    .din272_WIDTH( 16 ),
    .din273_WIDTH( 16 ),
    .din274_WIDTH( 16 ),
    .din275_WIDTH( 16 ),
    .din276_WIDTH( 16 ),
    .din277_WIDTH( 16 ),
    .din278_WIDTH( 16 ),
    .din279_WIDTH( 16 ),
    .din280_WIDTH( 16 ),
    .din281_WIDTH( 16 ),
    .din282_WIDTH( 16 ),
    .din283_WIDTH( 16 ),
    .din284_WIDTH( 16 ),
    .din285_WIDTH( 16 ),
    .din286_WIDTH( 16 ),
    .din287_WIDTH( 16 ),
    .din288_WIDTH( 16 ),
    .din289_WIDTH( 16 ),
    .din290_WIDTH( 16 ),
    .din291_WIDTH( 16 ),
    .din292_WIDTH( 16 ),
    .din293_WIDTH( 16 ),
    .din294_WIDTH( 16 ),
    .din295_WIDTH( 16 ),
    .din296_WIDTH( 16 ),
    .din297_WIDTH( 16 ),
    .din298_WIDTH( 16 ),
    .din299_WIDTH( 16 ),
    .din300_WIDTH( 16 ),
    .din301_WIDTH( 16 ),
    .din302_WIDTH( 16 ),
    .din303_WIDTH( 16 ),
    .din304_WIDTH( 16 ),
    .din305_WIDTH( 16 ),
    .din306_WIDTH( 16 ),
    .din307_WIDTH( 16 ),
    .din308_WIDTH( 16 ),
    .din309_WIDTH( 16 ),
    .din310_WIDTH( 16 ),
    .din311_WIDTH( 16 ),
    .din312_WIDTH( 16 ),
    .din313_WIDTH( 16 ),
    .din314_WIDTH( 16 ),
    .din315_WIDTH( 16 ),
    .din316_WIDTH( 16 ),
    .din317_WIDTH( 16 ),
    .din318_WIDTH( 16 ),
    .din319_WIDTH( 16 ),
    .din320_WIDTH( 16 ),
    .din321_WIDTH( 16 ),
    .din322_WIDTH( 16 ),
    .din323_WIDTH( 16 ),
    .din324_WIDTH( 16 ),
    .din325_WIDTH( 16 ),
    .din326_WIDTH( 16 ),
    .din327_WIDTH( 16 ),
    .din328_WIDTH( 16 ),
    .din329_WIDTH( 16 ),
    .din330_WIDTH( 16 ),
    .din331_WIDTH( 16 ),
    .din332_WIDTH( 16 ),
    .din333_WIDTH( 16 ),
    .din334_WIDTH( 16 ),
    .din335_WIDTH( 16 ),
    .din336_WIDTH( 16 ),
    .din337_WIDTH( 16 ),
    .din338_WIDTH( 16 ),
    .din339_WIDTH( 16 ),
    .din340_WIDTH( 16 ),
    .din341_WIDTH( 16 ),
    .din342_WIDTH( 16 ),
    .din343_WIDTH( 16 ),
    .din344_WIDTH( 16 ),
    .din345_WIDTH( 16 ),
    .din346_WIDTH( 16 ),
    .din347_WIDTH( 16 ),
    .din348_WIDTH( 16 ),
    .din349_WIDTH( 16 ),
    .din350_WIDTH( 16 ),
    .din351_WIDTH( 16 ),
    .din352_WIDTH( 16 ),
    .din353_WIDTH( 16 ),
    .din354_WIDTH( 16 ),
    .din355_WIDTH( 16 ),
    .din356_WIDTH( 16 ),
    .din357_WIDTH( 16 ),
    .din358_WIDTH( 16 ),
    .din359_WIDTH( 16 ),
    .din360_WIDTH( 16 ),
    .din361_WIDTH( 16 ),
    .din362_WIDTH( 16 ),
    .din363_WIDTH( 16 ),
    .din364_WIDTH( 16 ),
    .din365_WIDTH( 16 ),
    .din366_WIDTH( 16 ),
    .din367_WIDTH( 16 ),
    .din368_WIDTH( 16 ),
    .din369_WIDTH( 16 ),
    .din370_WIDTH( 16 ),
    .din371_WIDTH( 16 ),
    .din372_WIDTH( 16 ),
    .din373_WIDTH( 16 ),
    .din374_WIDTH( 16 ),
    .din375_WIDTH( 16 ),
    .din376_WIDTH( 16 ),
    .din377_WIDTH( 16 ),
    .din378_WIDTH( 16 ),
    .din379_WIDTH( 16 ),
    .din380_WIDTH( 16 ),
    .din381_WIDTH( 16 ),
    .din382_WIDTH( 16 ),
    .din383_WIDTH( 16 ),
    .din384_WIDTH( 16 ),
    .din385_WIDTH( 16 ),
    .din386_WIDTH( 16 ),
    .din387_WIDTH( 16 ),
    .din388_WIDTH( 16 ),
    .din389_WIDTH( 16 ),
    .din390_WIDTH( 16 ),
    .din391_WIDTH( 16 ),
    .din392_WIDTH( 16 ),
    .din393_WIDTH( 16 ),
    .din394_WIDTH( 16 ),
    .din395_WIDTH( 16 ),
    .din396_WIDTH( 16 ),
    .din397_WIDTH( 16 ),
    .din398_WIDTH( 16 ),
    .din399_WIDTH( 16 ),
    .din400_WIDTH( 16 ),
    .din401_WIDTH( 16 ),
    .din402_WIDTH( 16 ),
    .din403_WIDTH( 16 ),
    .din404_WIDTH( 16 ),
    .din405_WIDTH( 16 ),
    .din406_WIDTH( 16 ),
    .din407_WIDTH( 16 ),
    .din408_WIDTH( 16 ),
    .din409_WIDTH( 16 ),
    .din410_WIDTH( 16 ),
    .din411_WIDTH( 16 ),
    .din412_WIDTH( 16 ),
    .din413_WIDTH( 16 ),
    .din414_WIDTH( 16 ),
    .din415_WIDTH( 16 ),
    .din416_WIDTH( 16 ),
    .din417_WIDTH( 16 ),
    .din418_WIDTH( 16 ),
    .din419_WIDTH( 16 ),
    .din420_WIDTH( 16 ),
    .din421_WIDTH( 16 ),
    .din422_WIDTH( 16 ),
    .din423_WIDTH( 16 ),
    .din424_WIDTH( 16 ),
    .din425_WIDTH( 16 ),
    .din426_WIDTH( 16 ),
    .din427_WIDTH( 16 ),
    .din428_WIDTH( 16 ),
    .din429_WIDTH( 16 ),
    .din430_WIDTH( 16 ),
    .din431_WIDTH( 16 ),
    .din432_WIDTH( 16 ),
    .din433_WIDTH( 16 ),
    .din434_WIDTH( 16 ),
    .din435_WIDTH( 16 ),
    .din436_WIDTH( 16 ),
    .din437_WIDTH( 16 ),
    .din438_WIDTH( 16 ),
    .din439_WIDTH( 16 ),
    .din440_WIDTH( 16 ),
    .din441_WIDTH( 16 ),
    .din442_WIDTH( 16 ),
    .din443_WIDTH( 16 ),
    .din444_WIDTH( 16 ),
    .din445_WIDTH( 16 ),
    .din446_WIDTH( 16 ),
    .din447_WIDTH( 16 ),
    .din448_WIDTH( 16 ),
    .din449_WIDTH( 16 ),
    .din450_WIDTH( 16 ),
    .din451_WIDTH( 16 ),
    .din452_WIDTH( 16 ),
    .din453_WIDTH( 16 ),
    .din454_WIDTH( 16 ),
    .din455_WIDTH( 16 ),
    .din456_WIDTH( 16 ),
    .din457_WIDTH( 16 ),
    .din458_WIDTH( 16 ),
    .din459_WIDTH( 16 ),
    .din460_WIDTH( 16 ),
    .din461_WIDTH( 16 ),
    .din462_WIDTH( 16 ),
    .din463_WIDTH( 16 ),
    .din464_WIDTH( 16 ),
    .din465_WIDTH( 16 ),
    .din466_WIDTH( 16 ),
    .din467_WIDTH( 16 ),
    .din468_WIDTH( 16 ),
    .din469_WIDTH( 16 ),
    .din470_WIDTH( 16 ),
    .din471_WIDTH( 16 ),
    .din472_WIDTH( 16 ),
    .din473_WIDTH( 16 ),
    .din474_WIDTH( 16 ),
    .din475_WIDTH( 16 ),
    .din476_WIDTH( 16 ),
    .din477_WIDTH( 16 ),
    .din478_WIDTH( 16 ),
    .din479_WIDTH( 16 ),
    .din480_WIDTH( 16 ),
    .din481_WIDTH( 16 ),
    .din482_WIDTH( 16 ),
    .din483_WIDTH( 16 ),
    .din484_WIDTH( 16 ),
    .din485_WIDTH( 16 ),
    .din486_WIDTH( 16 ),
    .din487_WIDTH( 16 ),
    .din488_WIDTH( 16 ),
    .din489_WIDTH( 16 ),
    .din490_WIDTH( 16 ),
    .din491_WIDTH( 16 ),
    .din492_WIDTH( 16 ),
    .din493_WIDTH( 16 ),
    .din494_WIDTH( 16 ),
    .din495_WIDTH( 16 ),
    .din496_WIDTH( 16 ),
    .din497_WIDTH( 16 ),
    .din498_WIDTH( 16 ),
    .din499_WIDTH( 16 ),
    .din500_WIDTH( 16 ),
    .din501_WIDTH( 16 ),
    .din502_WIDTH( 16 ),
    .din503_WIDTH( 16 ),
    .din504_WIDTH( 16 ),
    .din505_WIDTH( 16 ),
    .din506_WIDTH( 16 ),
    .din507_WIDTH( 16 ),
    .din508_WIDTH( 16 ),
    .din509_WIDTH( 16 ),
    .din510_WIDTH( 16 ),
    .din511_WIDTH( 16 ),
    .din512_WIDTH( 16 ),
    .din513_WIDTH( 16 ),
    .din514_WIDTH( 16 ),
    .din515_WIDTH( 16 ),
    .din516_WIDTH( 16 ),
    .din517_WIDTH( 16 ),
    .din518_WIDTH( 16 ),
    .din519_WIDTH( 16 ),
    .din520_WIDTH( 16 ),
    .din521_WIDTH( 16 ),
    .din522_WIDTH( 16 ),
    .din523_WIDTH( 16 ),
    .din524_WIDTH( 16 ),
    .din525_WIDTH( 16 ),
    .din526_WIDTH( 16 ),
    .din527_WIDTH( 16 ),
    .din528_WIDTH( 16 ),
    .din529_WIDTH( 16 ),
    .din530_WIDTH( 16 ),
    .din531_WIDTH( 16 ),
    .din532_WIDTH( 16 ),
    .din533_WIDTH( 16 ),
    .din534_WIDTH( 16 ),
    .din535_WIDTH( 16 ),
    .din536_WIDTH( 16 ),
    .din537_WIDTH( 16 ),
    .din538_WIDTH( 16 ),
    .din539_WIDTH( 16 ),
    .din540_WIDTH( 16 ),
    .din541_WIDTH( 16 ),
    .din542_WIDTH( 16 ),
    .din543_WIDTH( 16 ),
    .din544_WIDTH( 16 ),
    .din545_WIDTH( 16 ),
    .din546_WIDTH( 16 ),
    .din547_WIDTH( 16 ),
    .din548_WIDTH( 16 ),
    .din549_WIDTH( 16 ),
    .din550_WIDTH( 16 ),
    .din551_WIDTH( 16 ),
    .din552_WIDTH( 16 ),
    .din553_WIDTH( 16 ),
    .din554_WIDTH( 16 ),
    .din555_WIDTH( 16 ),
    .din556_WIDTH( 16 ),
    .din557_WIDTH( 16 ),
    .din558_WIDTH( 16 ),
    .din559_WIDTH( 16 ),
    .din560_WIDTH( 16 ),
    .din561_WIDTH( 16 ),
    .din562_WIDTH( 16 ),
    .din563_WIDTH( 16 ),
    .din564_WIDTH( 16 ),
    .din565_WIDTH( 16 ),
    .din566_WIDTH( 16 ),
    .din567_WIDTH( 16 ),
    .din568_WIDTH( 16 ),
    .din569_WIDTH( 16 ),
    .din570_WIDTH( 16 ),
    .din571_WIDTH( 16 ),
    .din572_WIDTH( 16 ),
    .din573_WIDTH( 16 ),
    .din574_WIDTH( 16 ),
    .din575_WIDTH( 16 ),
    .din576_WIDTH( 10 ),
    .dout_WIDTH( 16 ))
StreamingFCLayer_5jm_U1(
    .din0(tmp_V_fu_1410),
    .din1(tmp_V_1_fu_1414),
    .din2(tmp_V_2_fu_1418),
    .din3(tmp_V_4_fu_1422),
    .din4(tmp_V_5_fu_1426),
    .din5(tmp_V_6_fu_1430),
    .din6(tmp_V_7_fu_1434),
    .din7(tmp_V_8_fu_1438),
    .din8(tmp_V_9_fu_1442),
    .din9(tmp_V_10_fu_1446),
    .din10(tmp_V_11_fu_1450),
    .din11(tmp_V_12_fu_1454),
    .din12(tmp_V_13_fu_1458),
    .din13(tmp_V_14_fu_1462),
    .din14(tmp_V_15_fu_1466),
    .din15(tmp_V_16_fu_1470),
    .din16(tmp_V_17_fu_1474),
    .din17(tmp_V_18_fu_1478),
    .din18(tmp_V_19_fu_1482),
    .din19(tmp_V_20_fu_1486),
    .din20(tmp_V_21_fu_1490),
    .din21(tmp_V_22_fu_1494),
    .din22(tmp_V_23_fu_1498),
    .din23(tmp_V_24_fu_1502),
    .din24(tmp_V_25_fu_1506),
    .din25(tmp_V_26_fu_1510),
    .din26(tmp_V_27_fu_1514),
    .din27(tmp_V_28_fu_1518),
    .din28(tmp_V_29_fu_1522),
    .din29(tmp_V_30_fu_1526),
    .din30(tmp_V_31_fu_1530),
    .din31(tmp_V_32_fu_1534),
    .din32(tmp_V_33_fu_1538),
    .din33(tmp_V_34_fu_1542),
    .din34(tmp_V_35_fu_1546),
    .din35(tmp_V_36_fu_1550),
    .din36(tmp_V_37_fu_1554),
    .din37(tmp_V_38_fu_1558),
    .din38(tmp_V_39_fu_1562),
    .din39(tmp_V_40_fu_1566),
    .din40(tmp_V_41_fu_1570),
    .din41(tmp_V_42_fu_1574),
    .din42(tmp_V_43_fu_1578),
    .din43(tmp_V_44_fu_1582),
    .din44(tmp_V_45_fu_1586),
    .din45(tmp_V_46_fu_1590),
    .din46(tmp_V_47_fu_1594),
    .din47(tmp_V_48_fu_1598),
    .din48(tmp_V_49_fu_1602),
    .din49(tmp_V_50_fu_1606),
    .din50(tmp_V_51_fu_1610),
    .din51(tmp_V_52_fu_1614),
    .din52(tmp_V_53_fu_1618),
    .din53(tmp_V_54_fu_1622),
    .din54(tmp_V_55_fu_1626),
    .din55(tmp_V_56_fu_1630),
    .din56(tmp_V_57_fu_1634),
    .din57(tmp_V_58_fu_1638),
    .din58(tmp_V_59_fu_1642),
    .din59(tmp_V_60_fu_1646),
    .din60(tmp_V_61_fu_1650),
    .din61(tmp_V_62_fu_1654),
    .din62(tmp_V_63_fu_1658),
    .din63(tmp_V_64_fu_1662),
    .din64(tmp_V_65_fu_1666),
    .din65(tmp_V_66_fu_1670),
    .din66(tmp_V_67_fu_1674),
    .din67(tmp_V_68_fu_1678),
    .din68(tmp_V_69_fu_1682),
    .din69(tmp_V_70_fu_1686),
    .din70(tmp_V_71_fu_1690),
    .din71(tmp_V_72_fu_1694),
    .din72(tmp_V_73_fu_1698),
    .din73(tmp_V_74_fu_1702),
    .din74(tmp_V_75_fu_1706),
    .din75(tmp_V_76_fu_1710),
    .din76(tmp_V_77_fu_1714),
    .din77(tmp_V_78_fu_1718),
    .din78(tmp_V_79_fu_1722),
    .din79(tmp_V_80_fu_1726),
    .din80(tmp_V_81_fu_1730),
    .din81(tmp_V_82_fu_1734),
    .din82(tmp_V_83_fu_1738),
    .din83(tmp_V_84_fu_1742),
    .din84(tmp_V_85_fu_1746),
    .din85(tmp_V_86_fu_1750),
    .din86(tmp_V_87_fu_1754),
    .din87(tmp_V_88_fu_1758),
    .din88(tmp_V_89_fu_1762),
    .din89(tmp_V_90_fu_1766),
    .din90(tmp_V_91_fu_1770),
    .din91(tmp_V_92_fu_1774),
    .din92(tmp_V_93_fu_1778),
    .din93(tmp_V_94_fu_1782),
    .din94(tmp_V_95_fu_1786),
    .din95(tmp_V_96_fu_1790),
    .din96(tmp_V_97_fu_1794),
    .din97(tmp_V_98_fu_1798),
    .din98(tmp_V_99_fu_1802),
    .din99(tmp_V_100_fu_1806),
    .din100(tmp_V_101_fu_1810),
    .din101(tmp_V_102_fu_1814),
    .din102(tmp_V_103_fu_1818),
    .din103(tmp_V_104_fu_1822),
    .din104(tmp_V_105_fu_1826),
    .din105(tmp_V_106_fu_1830),
    .din106(tmp_V_107_fu_1834),
    .din107(tmp_V_108_fu_1838),
    .din108(tmp_V_109_fu_1842),
    .din109(tmp_V_110_fu_1846),
    .din110(tmp_V_111_fu_1850),
    .din111(tmp_V_112_fu_1854),
    .din112(tmp_V_113_fu_1858),
    .din113(tmp_V_114_fu_1862),
    .din114(tmp_V_115_fu_1866),
    .din115(tmp_V_116_fu_1870),
    .din116(tmp_V_117_fu_1874),
    .din117(tmp_V_118_fu_1878),
    .din118(tmp_V_119_fu_1882),
    .din119(tmp_V_120_fu_1886),
    .din120(tmp_V_121_fu_1890),
    .din121(tmp_V_122_fu_1894),
    .din122(tmp_V_123_fu_1898),
    .din123(tmp_V_124_fu_1902),
    .din124(tmp_V_125_fu_1906),
    .din125(tmp_V_126_fu_1910),
    .din126(tmp_V_127_fu_1914),
    .din127(tmp_V_128_fu_1918),
    .din128(tmp_V_129_fu_1922),
    .din129(tmp_V_130_fu_1926),
    .din130(tmp_V_131_fu_1930),
    .din131(tmp_V_132_fu_1934),
    .din132(tmp_V_133_fu_1938),
    .din133(tmp_V_134_fu_1942),
    .din134(tmp_V_135_fu_1946),
    .din135(tmp_V_136_fu_1950),
    .din136(tmp_V_137_fu_1954),
    .din137(tmp_V_138_fu_1958),
    .din138(tmp_V_139_fu_1962),
    .din139(tmp_V_140_fu_1966),
    .din140(tmp_V_141_fu_1970),
    .din141(tmp_V_142_fu_1974),
    .din142(tmp_V_143_fu_1978),
    .din143(tmp_V_144_fu_1982),
    .din144(tmp_V_145_fu_1986),
    .din145(tmp_V_146_fu_1990),
    .din146(tmp_V_147_fu_1994),
    .din147(tmp_V_148_fu_1998),
    .din148(tmp_V_149_fu_2002),
    .din149(tmp_V_150_fu_2006),
    .din150(tmp_V_151_fu_2010),
    .din151(tmp_V_152_fu_2014),
    .din152(tmp_V_153_fu_2018),
    .din153(tmp_V_154_fu_2022),
    .din154(tmp_V_155_fu_2026),
    .din155(tmp_V_156_fu_2030),
    .din156(tmp_V_157_fu_2034),
    .din157(tmp_V_158_fu_2038),
    .din158(tmp_V_159_fu_2042),
    .din159(tmp_V_160_fu_2046),
    .din160(tmp_V_161_fu_2050),
    .din161(tmp_V_162_fu_2054),
    .din162(tmp_V_163_fu_2058),
    .din163(tmp_V_164_fu_2062),
    .din164(tmp_V_165_fu_2066),
    .din165(tmp_V_166_fu_2070),
    .din166(tmp_V_167_fu_2074),
    .din167(tmp_V_168_fu_2078),
    .din168(tmp_V_169_fu_2082),
    .din169(tmp_V_170_fu_2086),
    .din170(tmp_V_171_fu_2090),
    .din171(tmp_V_172_fu_2094),
    .din172(tmp_V_173_fu_2098),
    .din173(tmp_V_174_fu_2102),
    .din174(tmp_V_175_fu_2106),
    .din175(tmp_V_176_fu_2110),
    .din176(tmp_V_177_fu_2114),
    .din177(tmp_V_178_fu_2118),
    .din178(tmp_V_179_fu_2122),
    .din179(tmp_V_180_fu_2126),
    .din180(tmp_V_181_fu_2130),
    .din181(tmp_V_182_fu_2134),
    .din182(tmp_V_183_fu_2138),
    .din183(tmp_V_184_fu_2142),
    .din184(tmp_V_185_fu_2146),
    .din185(tmp_V_186_fu_2150),
    .din186(tmp_V_187_fu_2154),
    .din187(tmp_V_188_fu_2158),
    .din188(tmp_V_189_fu_2162),
    .din189(tmp_V_190_fu_2166),
    .din190(tmp_V_191_fu_2170),
    .din191(tmp_V_192_fu_2174),
    .din192(tmp_V_193_fu_2178),
    .din193(tmp_V_194_fu_2182),
    .din194(tmp_V_195_fu_2186),
    .din195(tmp_V_196_fu_2190),
    .din196(tmp_V_197_fu_2194),
    .din197(tmp_V_198_fu_2198),
    .din198(tmp_V_199_fu_2202),
    .din199(tmp_V_200_fu_2206),
    .din200(tmp_V_201_fu_2210),
    .din201(tmp_V_202_fu_2214),
    .din202(tmp_V_203_fu_2218),
    .din203(tmp_V_204_fu_2222),
    .din204(tmp_V_205_fu_2226),
    .din205(tmp_V_206_fu_2230),
    .din206(tmp_V_207_fu_2234),
    .din207(tmp_V_208_fu_2238),
    .din208(tmp_V_209_fu_2242),
    .din209(tmp_V_210_fu_2246),
    .din210(tmp_V_211_fu_2250),
    .din211(tmp_V_212_fu_2254),
    .din212(tmp_V_213_fu_2258),
    .din213(tmp_V_214_fu_2262),
    .din214(tmp_V_215_fu_2266),
    .din215(tmp_V_216_fu_2270),
    .din216(tmp_V_217_fu_2274),
    .din217(tmp_V_218_fu_2278),
    .din218(tmp_V_219_fu_2282),
    .din219(tmp_V_220_fu_2286),
    .din220(tmp_V_221_fu_2290),
    .din221(tmp_V_222_fu_2294),
    .din222(tmp_V_223_fu_2298),
    .din223(tmp_V_224_fu_2302),
    .din224(tmp_V_225_fu_2306),
    .din225(tmp_V_226_fu_2310),
    .din226(tmp_V_227_fu_2314),
    .din227(tmp_V_228_fu_2318),
    .din228(tmp_V_229_fu_2322),
    .din229(tmp_V_230_fu_2326),
    .din230(tmp_V_231_fu_2330),
    .din231(tmp_V_232_fu_2334),
    .din232(tmp_V_233_fu_2338),
    .din233(tmp_V_234_fu_2342),
    .din234(tmp_V_235_fu_2346),
    .din235(tmp_V_236_fu_2350),
    .din236(tmp_V_237_fu_2354),
    .din237(tmp_V_238_fu_2358),
    .din238(tmp_V_239_fu_2362),
    .din239(tmp_V_240_fu_2366),
    .din240(tmp_V_241_fu_2370),
    .din241(tmp_V_242_fu_2374),
    .din242(tmp_V_243_fu_2378),
    .din243(tmp_V_244_fu_2382),
    .din244(tmp_V_245_fu_2386),
    .din245(tmp_V_246_fu_2390),
    .din246(tmp_V_247_fu_2394),
    .din247(tmp_V_248_fu_2398),
    .din248(tmp_V_249_fu_2402),
    .din249(tmp_V_250_fu_2406),
    .din250(tmp_V_251_fu_2410),
    .din251(tmp_V_252_fu_2414),
    .din252(tmp_V_253_fu_2418),
    .din253(tmp_V_254_fu_2422),
    .din254(tmp_V_255_fu_2426),
    .din255(tmp_V_256_fu_2430),
    .din256(tmp_V_257_fu_2434),
    .din257(tmp_V_258_fu_2438),
    .din258(tmp_V_259_fu_2442),
    .din259(tmp_V_260_fu_2446),
    .din260(tmp_V_261_fu_2450),
    .din261(tmp_V_262_fu_2454),
    .din262(tmp_V_263_fu_2458),
    .din263(tmp_V_264_fu_2462),
    .din264(tmp_V_265_fu_2466),
    .din265(tmp_V_266_fu_2470),
    .din266(tmp_V_267_fu_2474),
    .din267(tmp_V_268_fu_2478),
    .din268(tmp_V_269_fu_2482),
    .din269(tmp_V_270_fu_2486),
    .din270(tmp_V_271_fu_2490),
    .din271(tmp_V_272_fu_2494),
    .din272(tmp_V_273_fu_2498),
    .din273(tmp_V_274_fu_2502),
    .din274(tmp_V_275_fu_2506),
    .din275(tmp_V_276_fu_2510),
    .din276(tmp_V_277_fu_2514),
    .din277(tmp_V_278_fu_2518),
    .din278(tmp_V_279_fu_2522),
    .din279(tmp_V_280_fu_2526),
    .din280(tmp_V_281_fu_2530),
    .din281(tmp_V_282_fu_2534),
    .din282(tmp_V_283_fu_2538),
    .din283(tmp_V_284_fu_2542),
    .din284(tmp_V_285_fu_2546),
    .din285(tmp_V_286_fu_2550),
    .din286(tmp_V_287_fu_2554),
    .din287(tmp_V_288_fu_2558),
    .din288(tmp_V_289_fu_2562),
    .din289(tmp_V_290_fu_2566),
    .din290(tmp_V_291_fu_2570),
    .din291(tmp_V_292_fu_2574),
    .din292(tmp_V_293_fu_2578),
    .din293(tmp_V_294_fu_2582),
    .din294(tmp_V_295_fu_2586),
    .din295(tmp_V_296_fu_2590),
    .din296(tmp_V_297_fu_2594),
    .din297(tmp_V_298_fu_2598),
    .din298(tmp_V_299_fu_2602),
    .din299(tmp_V_300_fu_2606),
    .din300(tmp_V_301_fu_2610),
    .din301(tmp_V_302_fu_2614),
    .din302(tmp_V_303_fu_2618),
    .din303(tmp_V_304_fu_2622),
    .din304(tmp_V_305_fu_2626),
    .din305(tmp_V_306_fu_2630),
    .din306(tmp_V_307_fu_2634),
    .din307(tmp_V_308_fu_2638),
    .din308(tmp_V_309_fu_2642),
    .din309(tmp_V_310_fu_2646),
    .din310(tmp_V_311_fu_2650),
    .din311(tmp_V_312_fu_2654),
    .din312(tmp_V_313_fu_2658),
    .din313(tmp_V_314_fu_2662),
    .din314(tmp_V_315_fu_2666),
    .din315(tmp_V_316_fu_2670),
    .din316(tmp_V_317_fu_2674),
    .din317(tmp_V_318_fu_2678),
    .din318(tmp_V_319_fu_2682),
    .din319(tmp_V_320_fu_2686),
    .din320(tmp_V_321_fu_2690),
    .din321(tmp_V_322_fu_2694),
    .din322(tmp_V_323_fu_2698),
    .din323(tmp_V_324_fu_2702),
    .din324(tmp_V_325_fu_2706),
    .din325(tmp_V_326_fu_2710),
    .din326(tmp_V_327_fu_2714),
    .din327(tmp_V_328_fu_2718),
    .din328(tmp_V_329_fu_2722),
    .din329(tmp_V_330_fu_2726),
    .din330(tmp_V_331_fu_2730),
    .din331(tmp_V_332_fu_2734),
    .din332(tmp_V_333_fu_2738),
    .din333(tmp_V_334_fu_2742),
    .din334(tmp_V_335_fu_2746),
    .din335(tmp_V_336_fu_2750),
    .din336(tmp_V_337_fu_2754),
    .din337(tmp_V_338_fu_2758),
    .din338(tmp_V_339_fu_2762),
    .din339(tmp_V_340_fu_2766),
    .din340(tmp_V_341_fu_2770),
    .din341(tmp_V_342_fu_2774),
    .din342(tmp_V_343_fu_2778),
    .din343(tmp_V_344_fu_2782),
    .din344(tmp_V_345_fu_2786),
    .din345(tmp_V_346_fu_2790),
    .din346(tmp_V_347_fu_2794),
    .din347(tmp_V_348_fu_2798),
    .din348(tmp_V_349_fu_2802),
    .din349(tmp_V_350_fu_2806),
    .din350(tmp_V_351_fu_2810),
    .din351(tmp_V_352_fu_2814),
    .din352(tmp_V_353_fu_2818),
    .din353(tmp_V_354_fu_2822),
    .din354(tmp_V_355_fu_2826),
    .din355(tmp_V_356_fu_2830),
    .din356(tmp_V_357_fu_2834),
    .din357(tmp_V_358_fu_2838),
    .din358(tmp_V_359_fu_2842),
    .din359(tmp_V_360_fu_2846),
    .din360(tmp_V_361_fu_2850),
    .din361(tmp_V_362_fu_2854),
    .din362(tmp_V_363_fu_2858),
    .din363(tmp_V_364_fu_2862),
    .din364(tmp_V_365_fu_2866),
    .din365(tmp_V_366_fu_2870),
    .din366(tmp_V_367_fu_2874),
    .din367(tmp_V_368_fu_2878),
    .din368(tmp_V_369_fu_2882),
    .din369(tmp_V_370_fu_2886),
    .din370(tmp_V_371_fu_2890),
    .din371(tmp_V_372_fu_2894),
    .din372(tmp_V_373_fu_2898),
    .din373(tmp_V_374_fu_2902),
    .din374(tmp_V_375_fu_2906),
    .din375(tmp_V_376_fu_2910),
    .din376(tmp_V_377_fu_2914),
    .din377(tmp_V_378_fu_2918),
    .din378(tmp_V_379_fu_2922),
    .din379(tmp_V_380_fu_2926),
    .din380(tmp_V_381_fu_2930),
    .din381(tmp_V_382_fu_2934),
    .din382(tmp_V_383_fu_2938),
    .din383(tmp_V_384_fu_2942),
    .din384(tmp_V_385_fu_2946),
    .din385(tmp_V_386_fu_2950),
    .din386(tmp_V_387_fu_2954),
    .din387(tmp_V_388_fu_2958),
    .din388(tmp_V_389_fu_2962),
    .din389(tmp_V_390_fu_2966),
    .din390(tmp_V_391_fu_2970),
    .din391(tmp_V_392_fu_2974),
    .din392(tmp_V_393_fu_2978),
    .din393(tmp_V_394_fu_2982),
    .din394(tmp_V_395_fu_2986),
    .din395(tmp_V_396_fu_2990),
    .din396(tmp_V_397_fu_2994),
    .din397(tmp_V_398_fu_2998),
    .din398(tmp_V_399_fu_3002),
    .din399(tmp_V_400_fu_3006),
    .din400(tmp_V_401_fu_3010),
    .din401(tmp_V_402_fu_3014),
    .din402(tmp_V_403_fu_3018),
    .din403(tmp_V_404_fu_3022),
    .din404(tmp_V_405_fu_3026),
    .din405(tmp_V_406_fu_3030),
    .din406(tmp_V_407_fu_3034),
    .din407(tmp_V_408_fu_3038),
    .din408(tmp_V_409_fu_3042),
    .din409(tmp_V_410_fu_3046),
    .din410(tmp_V_411_fu_3050),
    .din411(tmp_V_412_fu_3054),
    .din412(tmp_V_413_fu_3058),
    .din413(tmp_V_414_fu_3062),
    .din414(tmp_V_415_fu_3066),
    .din415(tmp_V_416_fu_3070),
    .din416(tmp_V_417_fu_3074),
    .din417(tmp_V_418_fu_3078),
    .din418(tmp_V_419_fu_3082),
    .din419(tmp_V_420_fu_3086),
    .din420(tmp_V_421_fu_3090),
    .din421(tmp_V_422_fu_3094),
    .din422(tmp_V_423_fu_3098),
    .din423(tmp_V_424_fu_3102),
    .din424(tmp_V_425_fu_3106),
    .din425(tmp_V_426_fu_3110),
    .din426(tmp_V_427_fu_3114),
    .din427(tmp_V_428_fu_3118),
    .din428(tmp_V_429_fu_3122),
    .din429(tmp_V_430_fu_3126),
    .din430(tmp_V_431_fu_3130),
    .din431(tmp_V_432_fu_3134),
    .din432(tmp_V_433_fu_3138),
    .din433(tmp_V_434_fu_3142),
    .din434(tmp_V_435_fu_3146),
    .din435(tmp_V_436_fu_3150),
    .din436(tmp_V_437_fu_3154),
    .din437(tmp_V_438_fu_3158),
    .din438(tmp_V_439_fu_3162),
    .din439(tmp_V_440_fu_3166),
    .din440(tmp_V_441_fu_3170),
    .din441(tmp_V_442_fu_3174),
    .din442(tmp_V_443_fu_3178),
    .din443(tmp_V_444_fu_3182),
    .din444(tmp_V_445_fu_3186),
    .din445(tmp_V_446_fu_3190),
    .din446(tmp_V_447_fu_3194),
    .din447(tmp_V_448_fu_3198),
    .din448(tmp_V_449_fu_3202),
    .din449(tmp_V_450_fu_3206),
    .din450(tmp_V_451_fu_3210),
    .din451(tmp_V_452_fu_3214),
    .din452(tmp_V_453_fu_3218),
    .din453(tmp_V_454_fu_3222),
    .din454(tmp_V_455_fu_3226),
    .din455(tmp_V_456_fu_3230),
    .din456(tmp_V_457_fu_3234),
    .din457(tmp_V_458_fu_3238),
    .din458(tmp_V_459_fu_3242),
    .din459(tmp_V_460_fu_3246),
    .din460(tmp_V_461_fu_3250),
    .din461(tmp_V_462_fu_3254),
    .din462(tmp_V_463_fu_3258),
    .din463(tmp_V_464_fu_3262),
    .din464(tmp_V_465_fu_3266),
    .din465(tmp_V_466_fu_3270),
    .din466(tmp_V_467_fu_3274),
    .din467(tmp_V_468_fu_3278),
    .din468(tmp_V_469_fu_3282),
    .din469(tmp_V_470_fu_3286),
    .din470(tmp_V_471_fu_3290),
    .din471(tmp_V_472_fu_3294),
    .din472(tmp_V_473_fu_3298),
    .din473(tmp_V_474_fu_3302),
    .din474(tmp_V_475_fu_3306),
    .din475(tmp_V_476_fu_3310),
    .din476(tmp_V_477_fu_3314),
    .din477(tmp_V_478_fu_3318),
    .din478(tmp_V_479_fu_3322),
    .din479(tmp_V_480_fu_3326),
    .din480(tmp_V_481_fu_3330),
    .din481(tmp_V_482_fu_3334),
    .din482(tmp_V_483_fu_3338),
    .din483(tmp_V_484_fu_3342),
    .din484(tmp_V_485_fu_3346),
    .din485(tmp_V_486_fu_3350),
    .din486(tmp_V_487_fu_3354),
    .din487(tmp_V_488_fu_3358),
    .din488(tmp_V_489_fu_3362),
    .din489(tmp_V_490_fu_3366),
    .din490(tmp_V_491_fu_3370),
    .din491(tmp_V_492_fu_3374),
    .din492(tmp_V_493_fu_3378),
    .din493(tmp_V_494_fu_3382),
    .din494(tmp_V_495_fu_3386),
    .din495(tmp_V_496_fu_3390),
    .din496(tmp_V_497_fu_3394),
    .din497(tmp_V_498_fu_3398),
    .din498(tmp_V_499_fu_3402),
    .din499(tmp_V_500_fu_3406),
    .din500(tmp_V_501_fu_3410),
    .din501(tmp_V_502_fu_3414),
    .din502(tmp_V_503_fu_3418),
    .din503(tmp_V_504_fu_3422),
    .din504(tmp_V_505_fu_3426),
    .din505(tmp_V_506_fu_3430),
    .din506(tmp_V_507_fu_3434),
    .din507(tmp_V_508_fu_3438),
    .din508(tmp_V_509_fu_3442),
    .din509(tmp_V_510_fu_3446),
    .din510(tmp_V_511_fu_3450),
    .din511(tmp_V_512_fu_3454),
    .din512(tmp_V_513_fu_3458),
    .din513(tmp_V_514_fu_3462),
    .din514(tmp_V_515_fu_3466),
    .din515(tmp_V_516_fu_3470),
    .din516(tmp_V_517_fu_3474),
    .din517(tmp_V_518_fu_3478),
    .din518(tmp_V_519_fu_3482),
    .din519(tmp_V_520_fu_3486),
    .din520(tmp_V_521_fu_3490),
    .din521(tmp_V_522_fu_3494),
    .din522(tmp_V_523_fu_3498),
    .din523(tmp_V_524_fu_3502),
    .din524(tmp_V_525_fu_3506),
    .din525(tmp_V_526_fu_3510),
    .din526(tmp_V_527_fu_3514),
    .din527(tmp_V_528_fu_3518),
    .din528(tmp_V_529_fu_3522),
    .din529(tmp_V_530_fu_3526),
    .din530(tmp_V_531_fu_3530),
    .din531(tmp_V_532_fu_3534),
    .din532(tmp_V_533_fu_3538),
    .din533(tmp_V_534_fu_3542),
    .din534(tmp_V_535_fu_3546),
    .din535(tmp_V_536_fu_3550),
    .din536(tmp_V_537_fu_3554),
    .din537(tmp_V_538_fu_3558),
    .din538(tmp_V_539_fu_3562),
    .din539(tmp_V_540_fu_3566),
    .din540(tmp_V_541_fu_3570),
    .din541(tmp_V_542_fu_3574),
    .din542(tmp_V_543_fu_3578),
    .din543(tmp_V_544_fu_3582),
    .din544(tmp_V_545_fu_3586),
    .din545(tmp_V_546_fu_3590),
    .din546(tmp_V_547_fu_3594),
    .din547(tmp_V_548_fu_3598),
    .din548(tmp_V_549_fu_3602),
    .din549(tmp_V_550_fu_3606),
    .din550(tmp_V_551_fu_3610),
    .din551(tmp_V_552_fu_3614),
    .din552(tmp_V_553_fu_3618),
    .din553(tmp_V_554_fu_3622),
    .din554(tmp_V_555_fu_3626),
    .din555(tmp_V_556_fu_3630),
    .din556(tmp_V_557_fu_3634),
    .din557(tmp_V_558_fu_3638),
    .din558(tmp_V_559_fu_3642),
    .din559(tmp_V_560_fu_3646),
    .din560(tmp_V_561_fu_3650),
    .din561(tmp_V_562_fu_3654),
    .din562(tmp_V_563_fu_3658),
    .din563(tmp_V_564_fu_3662),
    .din564(tmp_V_565_fu_3666),
    .din565(tmp_V_566_fu_3670),
    .din566(tmp_V_567_fu_3674),
    .din567(tmp_V_568_fu_3678),
    .din568(tmp_V_569_fu_3682),
    .din569(tmp_V_570_fu_3686),
    .din570(tmp_V_571_fu_3690),
    .din571(tmp_V_572_fu_3694),
    .din572(tmp_V_573_fu_3698),
    .din573(tmp_V_574_fu_3702),
    .din574(tmp_V_575_fu_3706),
    .din575(tmp_V_576_fu_3710),
    .din576(inElem_V_1_fu_7401_p577),
    .dout(inElem_V_1_fu_7401_p578)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U2(
    .din0(mul_ln1352_fu_11634_p0),
    .din1(trunc_ln647_reg_17688),
    .dout(mul_ln1352_fu_11634_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U3(
    .din0(mul_ln1352_1_fu_11661_p0),
    .din1(p_Result_1_0_1_reg_17693),
    .dout(mul_ln1352_1_fu_11661_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U4(
    .din0(mul_ln1352_2_fu_11684_p0),
    .din1(p_Result_1_0_2_reg_17698),
    .dout(mul_ln1352_2_fu_11684_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U5(
    .din0(mul_ln1352_3_fu_11711_p0),
    .din1(p_Result_1_0_3_reg_17703),
    .dout(mul_ln1352_3_fu_11711_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U6(
    .din0(mul_ln1352_4_fu_11736_p0),
    .din1(p_Result_1_1_reg_17708),
    .dout(mul_ln1352_4_fu_11736_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U7(
    .din0(mul_ln1352_5_fu_11749_p0),
    .din1(p_Result_1_1_1_reg_17713),
    .dout(mul_ln1352_5_fu_11749_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U8(
    .din0(mul_ln1352_6_fu_11758_p0),
    .din1(p_Result_1_1_2_reg_17718),
    .dout(mul_ln1352_6_fu_11758_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U9(
    .din0(mul_ln1352_7_fu_11771_p0),
    .din1(p_Result_1_1_3_reg_17723),
    .dout(mul_ln1352_7_fu_11771_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U10(
    .din0(mul_ln1352_8_fu_11796_p0),
    .din1(p_Result_1_2_reg_17728),
    .dout(mul_ln1352_8_fu_11796_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U11(
    .din0(mul_ln1352_9_fu_11809_p0),
    .din1(p_Result_1_2_1_reg_17733),
    .dout(mul_ln1352_9_fu_11809_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U12(
    .din0(mul_ln1352_10_fu_11818_p0),
    .din1(p_Result_1_2_2_reg_17738),
    .dout(mul_ln1352_10_fu_11818_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U13(
    .din0(mul_ln1352_11_fu_11831_p0),
    .din1(p_Result_1_2_3_reg_17743),
    .dout(mul_ln1352_11_fu_11831_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U14(
    .din0(mul_ln1352_12_fu_11856_p0),
    .din1(p_Result_1_3_reg_17748),
    .dout(mul_ln1352_12_fu_11856_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U15(
    .din0(mul_ln1352_13_fu_11869_p0),
    .din1(p_Result_1_3_1_reg_17753),
    .dout(mul_ln1352_13_fu_11869_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U16(
    .din0(mul_ln1352_14_fu_11878_p0),
    .din1(p_Result_1_3_2_reg_17758),
    .dout(mul_ln1352_14_fu_11878_p2)
);

StreamingFCLayer_Batch_1_StreamingFCLayer_6jw #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 4 ),
    .din1_WIDTH( 4 ),
    .dout_WIDTH( 8 ))
StreamingFCLayer_6jw_U17(
    .din0(mul_ln1352_15_fu_11891_p0),
    .din1(p_Result_1_3_3_reg_17763),
    .dout(mul_ln1352_15_fu_11891_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd0) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_4476 <= inElem_V_1_fu_7401_p578;
    end else if ((((trunc_ln321_fu_8559_p1 == 10'd46) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd45) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd44) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd43) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd42) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd41) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd40) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd39) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd38) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd37) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd36) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd35) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd34) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd33) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd32) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd31) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd30) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd29) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd28) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd27) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd26) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd25) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd24) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd23) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd22) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd21) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd20) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd19) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd18) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd17) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd16) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd15) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd14) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd13) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd12) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd11) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd10) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd9) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd8) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd7) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd6) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd5) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd4) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd3) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd2) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | (~(trunc_ln321_fu_8559_p1 == 10'd46) & ~(trunc_ln321_fu_8559_p1 == 10'd45) & ~(trunc_ln321_fu_8559_p1 == 10'd44) & ~(trunc_ln321_fu_8559_p1 == 10'd43) & ~(trunc_ln321_fu_8559_p1 == 10'd42) & ~(trunc_ln321_fu_8559_p1 == 10'd41) & ~(trunc_ln321_fu_8559_p1 == 10'd40) & ~(trunc_ln321_fu_8559_p1 == 10'd39) & ~(trunc_ln321_fu_8559_p1 == 10'd38) & ~(trunc_ln321_fu_8559_p1 == 10'd37) & ~(trunc_ln321_fu_8559_p1 == 10'd36) & ~(trunc_ln321_fu_8559_p1 == 10'd35) & ~(trunc_ln321_fu_8559_p1 == 10'd34) & ~(trunc_ln321_fu_8559_p1 == 10'd33) & ~(trunc_ln321_fu_8559_p1 == 10'd32) & ~(trunc_ln321_fu_8559_p1 == 10'd31) & ~(trunc_ln321_fu_8559_p1 == 10'd30) & ~(trunc_ln321_fu_8559_p1 == 10'd29) & ~(trunc_ln321_fu_8559_p1 == 10'd28) & ~(trunc_ln321_fu_8559_p1 == 10'd27) & ~(trunc_ln321_fu_8559_p1 == 10'd26) & ~(trunc_ln321_fu_8559_p1 == 10'd25) & ~(trunc_ln321_fu_8559_p1 == 10'd24) & ~(trunc_ln321_fu_8559_p1 == 10'd23) & ~(trunc_ln321_fu_8559_p1 == 10'd22) & ~(trunc_ln321_fu_8559_p1 == 10'd21) & ~(trunc_ln321_fu_8559_p1 == 10'd20) & ~(trunc_ln321_fu_8559_p1 == 10'd19) & ~(trunc_ln321_fu_8559_p1 == 10'd18) & ~(trunc_ln321_fu_8559_p1 == 10'd17) & ~(trunc_ln321_fu_8559_p1 == 10'd16) & ~(trunc_ln321_fu_8559_p1 == 10'd15) & ~(trunc_ln321_fu_8559_p1 == 10'd14) & ~(trunc_ln321_fu_8559_p1 == 10'd13) & ~(trunc_ln321_fu_8559_p1 == 10'd12) & ~(trunc_ln321_fu_8559_p1 == 10'd11) & ~(trunc_ln321_fu_8559_p1 == 10'd10) & ~(trunc_ln321_fu_8559_p1 == 10'd9) & ~(trunc_ln321_fu_8559_p1 == 10'd8) & ~(trunc_ln321_fu_8559_p1 == 10'd7) & ~(trunc_ln321_fu_8559_p1 == 10'd6) & ~(trunc_ln321_fu_8559_p1 == 10'd5) & ~(trunc_ln321_fu_8559_p1 == 10'd4) & ~(trunc_ln321_fu_8559_p1 == 10'd3) & ~(trunc_ln321_fu_8559_p1 == 10'd2) & ~(trunc_ln321_fu_8559_p1 == 10'd1) & ~(trunc_ln321_fu_8559_p1 == 10'd0) & ~(trunc_ln321_fu_8559_p1 == 10'd574) & ~(trunc_ln321_fu_8559_p1 == 10'd573) & ~(trunc_ln321_fu_8559_p1 == 10'd572) & ~(trunc_ln321_fu_8559_p1 == 10'd571) & ~(trunc_ln321_fu_8559_p1 == 10'd570) & ~(trunc_ln321_fu_8559_p1 == 10'd569) & ~(trunc_ln321_fu_8559_p1 == 10'd568) & ~(trunc_ln321_fu_8559_p1 == 10'd567) & ~(trunc_ln321_fu_8559_p1 == 10'd566) & ~(trunc_ln321_fu_8559_p1 == 10'd565) & ~(trunc_ln321_fu_8559_p1 == 10'd564) & ~(trunc_ln321_fu_8559_p1 == 10'd563) & ~(trunc_ln321_fu_8559_p1 == 10'd562) & ~(trunc_ln321_fu_8559_p1 == 10'd561) & ~(trunc_ln321_fu_8559_p1 == 10'd560) & ~(trunc_ln321_fu_8559_p1 == 10'd559) & ~(trunc_ln321_fu_8559_p1 == 10'd558) & ~(trunc_ln321_fu_8559_p1 == 10'd557) & ~(trunc_ln321_fu_8559_p1 == 10'd556) & ~(trunc_ln321_fu_8559_p1 == 10'd555) & ~(trunc_ln321_fu_8559_p1 == 10'd554) & ~(trunc_ln321_fu_8559_p1 == 10'd553) & ~(trunc_ln321_fu_8559_p1 == 10'd552) & ~(trunc_ln321_fu_8559_p1 == 10'd551) & ~(trunc_ln321_fu_8559_p1 == 10'd550) & ~(trunc_ln321_fu_8559_p1 == 10'd549) & ~(trunc_ln321_fu_8559_p1 == 10'd548) & ~(trunc_ln321_fu_8559_p1 == 10'd547) & ~(trunc_ln321_fu_8559_p1 == 10'd546) & ~(trunc_ln321_fu_8559_p1 == 10'd545) & ~(trunc_ln321_fu_8559_p1 == 10'd544) & ~(trunc_ln321_fu_8559_p1 == 10'd543) & ~(trunc_ln321_fu_8559_p1 == 10'd542) & ~(trunc_ln321_fu_8559_p1 == 10'd541) & ~(trunc_ln321_fu_8559_p1 == 10'd540) & ~(trunc_ln321_fu_8559_p1 == 10'd539) & ~(trunc_ln321_fu_8559_p1 == 10'd538) & ~(trunc_ln321_fu_8559_p1 == 10'd537) & ~(trunc_ln321_fu_8559_p1 == 10'd536) & ~(trunc_ln321_fu_8559_p1 == 10'd535) & ~(trunc_ln321_fu_8559_p1 == 10'd534) & ~(trunc_ln321_fu_8559_p1 == 10'd533) & ~(trunc_ln321_fu_8559_p1 == 10'd532) & ~(trunc_ln321_fu_8559_p1 == 10'd531) & ~(trunc_ln321_fu_8559_p1 == 10'd530) & ~(trunc_ln321_fu_8559_p1 == 10'd529) & ~(trunc_ln321_fu_8559_p1 == 10'd528) & ~(trunc_ln321_fu_8559_p1 == 10'd527) & ~(trunc_ln321_fu_8559_p1 == 10'd526) & ~(trunc_ln321_fu_8559_p1 == 10'd525) & ~(trunc_ln321_fu_8559_p1 == 10'd524) & ~(trunc_ln321_fu_8559_p1 == 10'd523) & ~(trunc_ln321_fu_8559_p1 == 10'd522) & ~(trunc_ln321_fu_8559_p1 == 10'd521) & ~(trunc_ln321_fu_8559_p1 == 10'd520) & ~(trunc_ln321_fu_8559_p1 == 10'd519) & ~(trunc_ln321_fu_8559_p1 == 10'd518) & ~(trunc_ln321_fu_8559_p1 == 10'd517) & ~(trunc_ln321_fu_8559_p1 == 10'd516) & ~(trunc_ln321_fu_8559_p1 == 10'd515) & ~(trunc_ln321_fu_8559_p1 == 10'd514) & ~(trunc_ln321_fu_8559_p1 == 10'd513) & ~(trunc_ln321_fu_8559_p1 == 10'd512) & ~(trunc_ln321_fu_8559_p1 == 10'd511) & ~(trunc_ln321_fu_8559_p1 == 10'd510) & ~(trunc_ln321_fu_8559_p1 == 10'd509) & ~(trunc_ln321_fu_8559_p1 == 10'd508) & ~(trunc_ln321_fu_8559_p1 == 10'd507) & ~(trunc_ln321_fu_8559_p1 == 10'd506) & ~(trunc_ln321_fu_8559_p1 == 10'd505) & ~(trunc_ln321_fu_8559_p1 == 10'd504) & ~(trunc_ln321_fu_8559_p1 == 10'd503) & ~(trunc_ln321_fu_8559_p1 == 10'd502) & ~(trunc_ln321_fu_8559_p1 == 10'd501) & ~(trunc_ln321_fu_8559_p1 == 10'd500) & ~(trunc_ln321_fu_8559_p1 == 10'd499) & ~(trunc_ln321_fu_8559_p1 == 10'd498) & ~(trunc_ln321_fu_8559_p1 == 10'd497) & ~(trunc_ln321_fu_8559_p1 == 10'd496) & ~(trunc_ln321_fu_8559_p1 == 10'd495) & ~(trunc_ln321_fu_8559_p1 == 10'd494) & ~(trunc_ln321_fu_8559_p1 == 10'd493) & ~(trunc_ln321_fu_8559_p1 == 10'd492) & ~(trunc_ln321_fu_8559_p1 == 10'd491) & ~(trunc_ln321_fu_8559_p1 == 10'd490) & ~(trunc_ln321_fu_8559_p1 == 10'd489) & ~(trunc_ln321_fu_8559_p1 == 10'd488) & ~(trunc_ln321_fu_8559_p1 == 10'd487) & ~(trunc_ln321_fu_8559_p1 == 10'd486) & ~(trunc_ln321_fu_8559_p1 == 10'd485) & ~(trunc_ln321_fu_8559_p1 == 10'd484) & ~(trunc_ln321_fu_8559_p1 == 10'd483) & ~(trunc_ln321_fu_8559_p1 == 10'd482) & ~(trunc_ln321_fu_8559_p1 == 10'd481) & ~(trunc_ln321_fu_8559_p1 == 10'd480) & ~(trunc_ln321_fu_8559_p1 == 10'd479) & ~(trunc_ln321_fu_8559_p1 == 10'd478) & ~(trunc_ln321_fu_8559_p1 == 10'd477) & ~(trunc_ln321_fu_8559_p1 == 10'd476) & ~(trunc_ln321_fu_8559_p1 == 10'd475) & ~(trunc_ln321_fu_8559_p1 == 10'd474) & ~(trunc_ln321_fu_8559_p1 == 10'd473) & ~(trunc_ln321_fu_8559_p1 == 10'd472) & ~(trunc_ln321_fu_8559_p1 == 10'd471) & ~(trunc_ln321_fu_8559_p1 == 10'd470) & ~(trunc_ln321_fu_8559_p1 == 10'd469) & ~(trunc_ln321_fu_8559_p1 == 10'd468) & ~(trunc_ln321_fu_8559_p1 == 10'd467) & ~(trunc_ln321_fu_8559_p1 == 10'd466) & ~(trunc_ln321_fu_8559_p1 == 10'd465) & ~(trunc_ln321_fu_8559_p1 == 10'd464) & ~(trunc_ln321_fu_8559_p1 == 10'd463) & ~(trunc_ln321_fu_8559_p1 == 10'd462) & ~(trunc_ln321_fu_8559_p1 == 10'd461) & ~(trunc_ln321_fu_8559_p1 == 10'd460) & ~(trunc_ln321_fu_8559_p1 == 10'd459) & ~(trunc_ln321_fu_8559_p1 == 10'd458) & ~(trunc_ln321_fu_8559_p1 == 10'd457) & ~(trunc_ln321_fu_8559_p1 == 10'd456) & ~(trunc_ln321_fu_8559_p1 == 10'd455) & ~(trunc_ln321_fu_8559_p1 == 10'd454) & ~(trunc_ln321_fu_8559_p1 == 10'd453) & ~(trunc_ln321_fu_8559_p1 == 10'd452) & ~(trunc_ln321_fu_8559_p1 == 10'd451) & ~(trunc_ln321_fu_8559_p1 == 10'd450) & ~(trunc_ln321_fu_8559_p1 == 10'd449) & ~(trunc_ln321_fu_8559_p1 == 10'd448) & ~(trunc_ln321_fu_8559_p1 == 10'd447) & ~(trunc_ln321_fu_8559_p1 == 10'd446) & ~(trunc_ln321_fu_8559_p1 == 10'd445) & ~(trunc_ln321_fu_8559_p1 == 10'd444) & ~(trunc_ln321_fu_8559_p1 == 10'd443) & ~(trunc_ln321_fu_8559_p1 == 10'd442) & ~(trunc_ln321_fu_8559_p1 == 10'd441) & ~(trunc_ln321_fu_8559_p1 == 10'd440) & ~(trunc_ln321_fu_8559_p1 == 10'd439) & ~(trunc_ln321_fu_8559_p1 == 10'd438) & ~(trunc_ln321_fu_8559_p1 == 10'd437) & ~(trunc_ln321_fu_8559_p1 == 10'd436) & ~(trunc_ln321_fu_8559_p1 == 10'd435) & ~(trunc_ln321_fu_8559_p1 == 10'd434) & ~(trunc_ln321_fu_8559_p1 == 10'd433) & ~(trunc_ln321_fu_8559_p1 == 10'd432) & ~(trunc_ln321_fu_8559_p1 == 10'd431) & ~(trunc_ln321_fu_8559_p1 == 10'd430) & ~(trunc_ln321_fu_8559_p1 == 10'd429) & ~(trunc_ln321_fu_8559_p1 == 10'd428) & ~(trunc_ln321_fu_8559_p1 == 10'd427) & ~(trunc_ln321_fu_8559_p1 == 10'd426) & ~(trunc_ln321_fu_8559_p1 == 10'd425) & ~(trunc_ln321_fu_8559_p1 == 10'd424) & ~(trunc_ln321_fu_8559_p1 == 10'd423) & ~(trunc_ln321_fu_8559_p1 == 10'd422) & ~(trunc_ln321_fu_8559_p1 == 10'd421) & ~(trunc_ln321_fu_8559_p1 == 10'd420) & ~(trunc_ln321_fu_8559_p1 == 10'd419) & ~(trunc_ln321_fu_8559_p1 == 10'd418) & ~(trunc_ln321_fu_8559_p1 == 10'd417) & ~(trunc_ln321_fu_8559_p1 == 10'd416) & ~(trunc_ln321_fu_8559_p1 == 10'd415) & ~(trunc_ln321_fu_8559_p1 == 10'd414) & ~(trunc_ln321_fu_8559_p1 == 10'd413) & ~(trunc_ln321_fu_8559_p1 == 10'd412) & ~(trunc_ln321_fu_8559_p1 == 10'd411) & ~(trunc_ln321_fu_8559_p1 == 10'd410) & ~(trunc_ln321_fu_8559_p1 == 10'd409) & ~(trunc_ln321_fu_8559_p1 == 10'd408) & ~(trunc_ln321_fu_8559_p1 == 10'd407) & ~(trunc_ln321_fu_8559_p1 == 10'd406) & ~(trunc_ln321_fu_8559_p1 == 10'd405) & ~(trunc_ln321_fu_8559_p1 == 10'd404) & ~(trunc_ln321_fu_8559_p1 == 10'd403) & ~(trunc_ln321_fu_8559_p1 == 10'd402) & ~(trunc_ln321_fu_8559_p1 == 10'd401) & ~(trunc_ln321_fu_8559_p1 == 10'd400) & ~(trunc_ln321_fu_8559_p1 == 10'd399) & ~(trunc_ln321_fu_8559_p1 == 10'd398) & ~(trunc_ln321_fu_8559_p1 == 10'd397) & ~(trunc_ln321_fu_8559_p1 == 10'd396) & ~(trunc_ln321_fu_8559_p1 == 10'd395) & ~(trunc_ln321_fu_8559_p1 == 10'd394) & ~(trunc_ln321_fu_8559_p1 == 10'd393) & ~(trunc_ln321_fu_8559_p1 == 10'd392) & ~(trunc_ln321_fu_8559_p1 == 10'd391) & ~(trunc_ln321_fu_8559_p1 == 10'd390) & ~(trunc_ln321_fu_8559_p1 == 10'd389) & ~(trunc_ln321_fu_8559_p1 == 10'd388) & ~(trunc_ln321_fu_8559_p1 == 10'd387) & ~(trunc_ln321_fu_8559_p1 == 10'd386) & ~(trunc_ln321_fu_8559_p1 == 10'd385) & ~(trunc_ln321_fu_8559_p1 == 10'd384) & ~(trunc_ln321_fu_8559_p1 == 10'd383) & ~(trunc_ln321_fu_8559_p1 == 10'd382) & ~(trunc_ln321_fu_8559_p1 == 10'd381) & ~(trunc_ln321_fu_8559_p1 == 10'd380) & ~(trunc_ln321_fu_8559_p1 == 10'd379) & ~(trunc_ln321_fu_8559_p1 == 10'd378) & ~(trunc_ln321_fu_8559_p1 == 10'd377) & ~(trunc_ln321_fu_8559_p1 == 10'd376) & ~(trunc_ln321_fu_8559_p1 == 10'd375) & ~(trunc_ln321_fu_8559_p1 == 10'd374) & ~(trunc_ln321_fu_8559_p1 == 10'd373) & ~(trunc_ln321_fu_8559_p1 == 10'd372) & ~(trunc_ln321_fu_8559_p1 == 10'd371) & ~(trunc_ln321_fu_8559_p1 == 10'd370) & ~(trunc_ln321_fu_8559_p1 == 10'd369) & ~(trunc_ln321_fu_8559_p1 == 10'd368) & ~(trunc_ln321_fu_8559_p1 == 10'd367) & ~(trunc_ln321_fu_8559_p1 == 10'd366) & ~(trunc_ln321_fu_8559_p1 == 10'd365) & ~(trunc_ln321_fu_8559_p1 == 10'd364) & ~(trunc_ln321_fu_8559_p1 == 10'd363) & ~(trunc_ln321_fu_8559_p1 == 10'd362) & ~(trunc_ln321_fu_8559_p1 == 10'd361) & ~(trunc_ln321_fu_8559_p1 == 10'd360) & ~(trunc_ln321_fu_8559_p1 == 10'd359) & ~(trunc_ln321_fu_8559_p1 == 10'd358) & ~(trunc_ln321_fu_8559_p1 == 10'd357) & ~(trunc_ln321_fu_8559_p1 == 10'd356) & ~(trunc_ln321_fu_8559_p1 == 10'd355) & ~(trunc_ln321_fu_8559_p1 == 10'd354) & ~(trunc_ln321_fu_8559_p1 == 10'd353) & ~(trunc_ln321_fu_8559_p1 == 10'd352) & ~(trunc_ln321_fu_8559_p1 == 10'd351) & ~(trunc_ln321_fu_8559_p1 == 10'd350) & ~(trunc_ln321_fu_8559_p1 == 10'd349) & ~(trunc_ln321_fu_8559_p1 == 10'd348) & ~(trunc_ln321_fu_8559_p1 == 10'd347) & ~(trunc_ln321_fu_8559_p1 == 10'd346) & ~(trunc_ln321_fu_8559_p1 == 10'd345) & ~(trunc_ln321_fu_8559_p1 == 10'd344) & ~(trunc_ln321_fu_8559_p1 == 10'd343) & ~(trunc_ln321_fu_8559_p1 == 10'd342) & ~(trunc_ln321_fu_8559_p1 == 10'd341) & ~(trunc_ln321_fu_8559_p1 == 10'd340) & ~(trunc_ln321_fu_8559_p1 == 10'd339) & ~(trunc_ln321_fu_8559_p1 == 10'd338) & ~(trunc_ln321_fu_8559_p1 == 10'd337) & ~(trunc_ln321_fu_8559_p1 == 10'd336) & ~(trunc_ln321_fu_8559_p1 == 10'd335) & ~(trunc_ln321_fu_8559_p1 == 10'd334) & ~(trunc_ln321_fu_8559_p1 == 10'd333) & ~(trunc_ln321_fu_8559_p1 == 10'd332) & ~(trunc_ln321_fu_8559_p1 == 10'd331) & ~(trunc_ln321_fu_8559_p1 == 10'd330) & ~(trunc_ln321_fu_8559_p1 == 10'd329) & ~(trunc_ln321_fu_8559_p1 == 10'd328) & ~(trunc_ln321_fu_8559_p1 == 10'd327) & ~(trunc_ln321_fu_8559_p1 == 10'd326) & ~(trunc_ln321_fu_8559_p1 == 10'd325) & ~(trunc_ln321_fu_8559_p1 == 10'd324) & ~(trunc_ln321_fu_8559_p1 == 10'd323) & ~(trunc_ln321_fu_8559_p1 == 10'd322) & ~(trunc_ln321_fu_8559_p1 == 10'd321) & ~(trunc_ln321_fu_8559_p1 == 10'd320) & ~(trunc_ln321_fu_8559_p1 == 10'd319) & ~(trunc_ln321_fu_8559_p1 == 10'd318) & ~(trunc_ln321_fu_8559_p1 == 10'd317) & ~(trunc_ln321_fu_8559_p1 == 10'd316) & ~(trunc_ln321_fu_8559_p1 == 10'd315) & ~(trunc_ln321_fu_8559_p1 == 10'd314) & ~(trunc_ln321_fu_8559_p1 == 10'd313) & ~(trunc_ln321_fu_8559_p1 == 10'd312) & ~(trunc_ln321_fu_8559_p1 == 10'd311) & ~(trunc_ln321_fu_8559_p1 == 10'd310) & ~(trunc_ln321_fu_8559_p1 == 10'd309) & ~(trunc_ln321_fu_8559_p1 == 10'd308) & ~(trunc_ln321_fu_8559_p1 == 10'd307) & ~(trunc_ln321_fu_8559_p1 == 10'd306) & ~(trunc_ln321_fu_8559_p1 == 10'd305) & ~(trunc_ln321_fu_8559_p1 == 10'd304) & ~(trunc_ln321_fu_8559_p1 == 10'd303) & ~(trunc_ln321_fu_8559_p1 == 10'd302) & ~(trunc_ln321_fu_8559_p1 == 10'd301) & ~(trunc_ln321_fu_8559_p1 == 10'd300) & ~(trunc_ln321_fu_8559_p1 == 10'd299) & ~(trunc_ln321_fu_8559_p1 == 10'd298) & ~(trunc_ln321_fu_8559_p1 == 10'd297) & ~(trunc_ln321_fu_8559_p1 == 10'd296) & ~(trunc_ln321_fu_8559_p1 == 10'd295) & ~(trunc_ln321_fu_8559_p1 == 10'd294) & ~(trunc_ln321_fu_8559_p1 == 10'd293) & ~(trunc_ln321_fu_8559_p1 == 10'd292) & ~(trunc_ln321_fu_8559_p1 == 10'd291) & ~(trunc_ln321_fu_8559_p1 == 10'd290) & ~(trunc_ln321_fu_8559_p1 == 10'd289) & ~(trunc_ln321_fu_8559_p1 == 10'd288) & ~(trunc_ln321_fu_8559_p1 == 10'd287) & ~(trunc_ln321_fu_8559_p1 == 10'd286) & ~(trunc_ln321_fu_8559_p1 == 10'd285) & ~(trunc_ln321_fu_8559_p1 == 10'd284) & ~(trunc_ln321_fu_8559_p1 == 10'd283) & ~(trunc_ln321_fu_8559_p1 == 10'd282) & ~(trunc_ln321_fu_8559_p1 == 10'd281) & ~(trunc_ln321_fu_8559_p1 == 10'd280) & ~(trunc_ln321_fu_8559_p1 == 10'd279) & ~(trunc_ln321_fu_8559_p1 == 10'd278) & ~(trunc_ln321_fu_8559_p1 == 10'd277) & ~(trunc_ln321_fu_8559_p1 == 10'd276) & ~(trunc_ln321_fu_8559_p1 == 10'd275) & ~(trunc_ln321_fu_8559_p1 == 10'd274) & ~(trunc_ln321_fu_8559_p1 == 10'd273) & ~(trunc_ln321_fu_8559_p1 == 10'd272) & ~(trunc_ln321_fu_8559_p1 == 10'd271) & ~(trunc_ln321_fu_8559_p1 == 10'd270) & ~(trunc_ln321_fu_8559_p1 == 10'd269) & ~(trunc_ln321_fu_8559_p1 == 10'd268) & ~(trunc_ln321_fu_8559_p1 == 10'd267) & ~(trunc_ln321_fu_8559_p1 == 10'd266) & ~(trunc_ln321_fu_8559_p1 == 10'd265) & ~(trunc_ln321_fu_8559_p1 == 10'd264) & ~(trunc_ln321_fu_8559_p1 == 10'd263) & ~(trunc_ln321_fu_8559_p1 == 10'd262) & ~(trunc_ln321_fu_8559_p1 == 10'd261) & ~(trunc_ln321_fu_8559_p1 == 10'd260) & ~(trunc_ln321_fu_8559_p1 == 10'd259) & ~(trunc_ln321_fu_8559_p1 == 10'd258) & ~(trunc_ln321_fu_8559_p1 == 10'd257) & ~(trunc_ln321_fu_8559_p1 == 10'd256) & ~(trunc_ln321_fu_8559_p1 == 10'd255) & ~(trunc_ln321_fu_8559_p1 == 10'd254) & ~(trunc_ln321_fu_8559_p1 == 10'd253) & ~(trunc_ln321_fu_8559_p1 == 10'd252) & ~(trunc_ln321_fu_8559_p1 == 10'd251) & ~(trunc_ln321_fu_8559_p1 == 10'd250) & ~(trunc_ln321_fu_8559_p1 == 10'd249) & ~(trunc_ln321_fu_8559_p1 == 10'd248) & ~(trunc_ln321_fu_8559_p1 == 10'd247) & ~(trunc_ln321_fu_8559_p1 == 10'd246) & ~(trunc_ln321_fu_8559_p1 == 10'd245) & ~(trunc_ln321_fu_8559_p1 == 10'd244) & ~(trunc_ln321_fu_8559_p1 == 10'd243) & ~(trunc_ln321_fu_8559_p1 == 10'd242) & ~(trunc_ln321_fu_8559_p1 == 10'd241) & ~(trunc_ln321_fu_8559_p1 == 10'd240) & ~(trunc_ln321_fu_8559_p1 == 10'd239) & ~(trunc_ln321_fu_8559_p1 == 10'd238) & ~(trunc_ln321_fu_8559_p1 == 10'd237) & ~(trunc_ln321_fu_8559_p1 == 10'd236) & ~(trunc_ln321_fu_8559_p1 == 10'd235) & ~(trunc_ln321_fu_8559_p1 == 10'd234) & ~(trunc_ln321_fu_8559_p1 == 10'd233) & ~(trunc_ln321_fu_8559_p1 == 10'd232) & ~(trunc_ln321_fu_8559_p1 == 10'd231) & ~(trunc_ln321_fu_8559_p1 == 10'd230) & ~(trunc_ln321_fu_8559_p1 == 10'd229) & ~(trunc_ln321_fu_8559_p1 == 10'd228) & ~(trunc_ln321_fu_8559_p1 == 10'd227) & ~(trunc_ln321_fu_8559_p1 == 10'd226) & ~(trunc_ln321_fu_8559_p1 == 10'd225) & ~(trunc_ln321_fu_8559_p1 == 10'd224) & ~(trunc_ln321_fu_8559_p1 == 10'd223) & ~(trunc_ln321_fu_8559_p1 == 10'd222) & ~(trunc_ln321_fu_8559_p1 == 10'd221) & ~(trunc_ln321_fu_8559_p1 == 10'd220) & ~(trunc_ln321_fu_8559_p1 == 10'd219) & ~(trunc_ln321_fu_8559_p1 == 10'd218) & ~(trunc_ln321_fu_8559_p1 == 10'd217) & ~(trunc_ln321_fu_8559_p1 == 10'd216) & ~(trunc_ln321_fu_8559_p1 == 10'd215) & ~(trunc_ln321_fu_8559_p1 == 10'd214) & ~(trunc_ln321_fu_8559_p1 == 10'd213) & ~(trunc_ln321_fu_8559_p1 == 10'd212) & ~(trunc_ln321_fu_8559_p1 == 10'd211) & ~(trunc_ln321_fu_8559_p1 == 10'd210) & ~(trunc_ln321_fu_8559_p1 == 10'd209) & ~(trunc_ln321_fu_8559_p1 == 10'd208) & ~(trunc_ln321_fu_8559_p1 == 10'd207) & ~(trunc_ln321_fu_8559_p1 == 10'd206) & ~(trunc_ln321_fu_8559_p1 == 10'd205) & ~(trunc_ln321_fu_8559_p1 == 10'd204) & ~(trunc_ln321_fu_8559_p1 == 10'd203) & ~(trunc_ln321_fu_8559_p1 == 10'd202) & ~(trunc_ln321_fu_8559_p1 == 10'd201) & ~(trunc_ln321_fu_8559_p1 == 10'd200) & ~(trunc_ln321_fu_8559_p1 == 10'd199) & ~(trunc_ln321_fu_8559_p1 == 10'd198) & ~(trunc_ln321_fu_8559_p1 == 10'd197) & ~(trunc_ln321_fu_8559_p1 == 10'd196) & ~(trunc_ln321_fu_8559_p1 == 10'd195) & ~(trunc_ln321_fu_8559_p1 == 10'd194) & ~(trunc_ln321_fu_8559_p1 == 10'd193) & ~(trunc_ln321_fu_8559_p1 == 10'd192) & ~(trunc_ln321_fu_8559_p1 == 10'd191) & ~(trunc_ln321_fu_8559_p1 == 10'd190) & ~(trunc_ln321_fu_8559_p1 == 10'd189) & ~(trunc_ln321_fu_8559_p1 == 10'd188) & ~(trunc_ln321_fu_8559_p1 == 10'd187) & ~(trunc_ln321_fu_8559_p1 == 10'd186) & ~(trunc_ln321_fu_8559_p1 == 10'd185) & ~(trunc_ln321_fu_8559_p1 == 10'd184) & ~(trunc_ln321_fu_8559_p1 == 10'd183) & ~(trunc_ln321_fu_8559_p1 == 10'd182) & ~(trunc_ln321_fu_8559_p1 == 10'd181) & ~(trunc_ln321_fu_8559_p1 == 10'd180) & ~(trunc_ln321_fu_8559_p1 == 10'd179) & ~(trunc_ln321_fu_8559_p1 == 10'd178) & ~(trunc_ln321_fu_8559_p1 == 10'd177) & ~(trunc_ln321_fu_8559_p1 == 10'd176) & ~(trunc_ln321_fu_8559_p1 == 10'd175) & ~(trunc_ln321_fu_8559_p1 == 10'd174) & ~(trunc_ln321_fu_8559_p1 == 10'd173) & ~(trunc_ln321_fu_8559_p1 == 10'd172) & ~(trunc_ln321_fu_8559_p1 == 10'd171) & ~(trunc_ln321_fu_8559_p1 == 10'd170) & ~(trunc_ln321_fu_8559_p1 == 10'd169) & ~(trunc_ln321_fu_8559_p1 == 10'd168) & ~(trunc_ln321_fu_8559_p1 == 10'd167) & ~(trunc_ln321_fu_8559_p1 == 10'd166) & ~(trunc_ln321_fu_8559_p1 == 10'd165) & ~(trunc_ln321_fu_8559_p1 == 10'd164) & ~(trunc_ln321_fu_8559_p1 == 10'd163) & ~(trunc_ln321_fu_8559_p1 == 10'd162) & ~(trunc_ln321_fu_8559_p1 == 10'd161) & ~(trunc_ln321_fu_8559_p1 == 10'd160) & ~(trunc_ln321_fu_8559_p1 == 10'd159) & ~(trunc_ln321_fu_8559_p1 == 10'd158) & ~(trunc_ln321_fu_8559_p1 == 10'd157) & ~(trunc_ln321_fu_8559_p1 == 10'd156) & ~(trunc_ln321_fu_8559_p1 == 10'd155) & ~(trunc_ln321_fu_8559_p1 == 10'd154) & ~(trunc_ln321_fu_8559_p1 == 10'd153) & ~(trunc_ln321_fu_8559_p1 == 10'd152) & ~(trunc_ln321_fu_8559_p1 == 10'd151) & ~(trunc_ln321_fu_8559_p1 == 10'd150) & ~(trunc_ln321_fu_8559_p1 == 10'd149) & ~(trunc_ln321_fu_8559_p1 == 10'd148) & ~(trunc_ln321_fu_8559_p1 == 10'd147) & ~(trunc_ln321_fu_8559_p1 == 10'd146) & ~(trunc_ln321_fu_8559_p1 == 10'd145) & ~(trunc_ln321_fu_8559_p1 == 10'd144) & ~(trunc_ln321_fu_8559_p1 == 10'd143) & ~(trunc_ln321_fu_8559_p1 == 10'd142) & ~(trunc_ln321_fu_8559_p1 == 10'd141) & ~(trunc_ln321_fu_8559_p1 == 10'd140) & ~(trunc_ln321_fu_8559_p1 == 10'd139) & ~(trunc_ln321_fu_8559_p1 == 10'd138) & ~(trunc_ln321_fu_8559_p1 == 10'd137) & ~(trunc_ln321_fu_8559_p1 == 10'd136) & ~(trunc_ln321_fu_8559_p1 == 10'd135) & ~(trunc_ln321_fu_8559_p1 == 10'd134) & ~(trunc_ln321_fu_8559_p1 == 10'd133) & ~(trunc_ln321_fu_8559_p1 == 10'd132) & ~(trunc_ln321_fu_8559_p1 == 10'd131) & ~(trunc_ln321_fu_8559_p1 == 10'd130) & ~(trunc_ln321_fu_8559_p1 == 10'd129) & ~(trunc_ln321_fu_8559_p1 == 10'd128) & ~(trunc_ln321_fu_8559_p1 == 10'd127) & ~(trunc_ln321_fu_8559_p1 == 10'd126) & ~(trunc_ln321_fu_8559_p1 == 10'd125) & ~(trunc_ln321_fu_8559_p1 == 10'd124) & ~(trunc_ln321_fu_8559_p1 == 10'd123) & ~(trunc_ln321_fu_8559_p1 == 10'd122) & ~(trunc_ln321_fu_8559_p1 == 10'd121) & ~(trunc_ln321_fu_8559_p1 == 10'd120) & ~(trunc_ln321_fu_8559_p1 == 10'd119) & ~(trunc_ln321_fu_8559_p1 == 10'd118) & ~(trunc_ln321_fu_8559_p1 == 10'd117) & ~(trunc_ln321_fu_8559_p1 == 10'd116) & ~(trunc_ln321_fu_8559_p1 == 10'd115) & ~(trunc_ln321_fu_8559_p1 == 10'd114) & ~(trunc_ln321_fu_8559_p1 == 10'd113) & ~(trunc_ln321_fu_8559_p1 == 10'd112) & ~(trunc_ln321_fu_8559_p1 == 10'd111) & ~(trunc_ln321_fu_8559_p1 == 10'd110) & ~(trunc_ln321_fu_8559_p1 == 10'd109) & ~(trunc_ln321_fu_8559_p1 == 10'd108) & ~(trunc_ln321_fu_8559_p1 == 10'd107) & ~(trunc_ln321_fu_8559_p1 == 10'd106) & ~(trunc_ln321_fu_8559_p1 == 10'd105) & ~(trunc_ln321_fu_8559_p1 == 10'd104) & ~(trunc_ln321_fu_8559_p1 == 10'd103) & ~(trunc_ln321_fu_8559_p1 == 10'd102) & ~(trunc_ln321_fu_8559_p1 == 10'd101) & ~(trunc_ln321_fu_8559_p1 == 10'd100) & ~(trunc_ln321_fu_8559_p1 == 10'd99) & ~(trunc_ln321_fu_8559_p1 == 10'd98) & ~(trunc_ln321_fu_8559_p1 == 10'd97) & ~(trunc_ln321_fu_8559_p1 == 10'd96) & ~(trunc_ln321_fu_8559_p1 == 10'd95) & ~(trunc_ln321_fu_8559_p1 == 10'd94) & ~(trunc_ln321_fu_8559_p1 == 10'd93) & ~(trunc_ln321_fu_8559_p1 == 10'd92) & ~(trunc_ln321_fu_8559_p1 == 10'd91) & ~(trunc_ln321_fu_8559_p1 == 10'd90) & ~(trunc_ln321_fu_8559_p1 == 10'd89) & ~(trunc_ln321_fu_8559_p1 == 10'd88) & ~(trunc_ln321_fu_8559_p1 == 10'd87) & ~(trunc_ln321_fu_8559_p1 == 10'd86) & ~(trunc_ln321_fu_8559_p1 == 10'd85) & ~(trunc_ln321_fu_8559_p1 == 10'd84) & ~(trunc_ln321_fu_8559_p1 == 10'd83) & ~(trunc_ln321_fu_8559_p1 == 10'd82) & ~(trunc_ln321_fu_8559_p1 == 10'd81) & ~(trunc_ln321_fu_8559_p1 == 10'd80) & ~(trunc_ln321_fu_8559_p1 == 10'd79) & ~(trunc_ln321_fu_8559_p1 == 10'd78) & ~(trunc_ln321_fu_8559_p1 == 10'd77) & ~(trunc_ln321_fu_8559_p1 == 10'd76) & ~(trunc_ln321_fu_8559_p1 == 10'd75) & ~(trunc_ln321_fu_8559_p1 == 10'd74) & ~(trunc_ln321_fu_8559_p1 == 10'd73) & ~(trunc_ln321_fu_8559_p1 == 10'd72) & ~(trunc_ln321_fu_8559_p1 == 10'd71) & ~(trunc_ln321_fu_8559_p1 == 10'd70) & ~(trunc_ln321_fu_8559_p1 == 10'd69) & ~(trunc_ln321_fu_8559_p1 == 10'd68) & ~(trunc_ln321_fu_8559_p1 == 10'd67) & ~(trunc_ln321_fu_8559_p1 == 10'd66) & ~(trunc_ln321_fu_8559_p1 == 10'd65) & ~(trunc_ln321_fu_8559_p1 == 10'd64) & ~(trunc_ln321_fu_8559_p1 == 10'd63) & ~(trunc_ln321_fu_8559_p1 == 10'd62) & ~(trunc_ln321_fu_8559_p1 == 10'd61) & ~(trunc_ln321_fu_8559_p1 == 10'd60) & ~(trunc_ln321_fu_8559_p1 == 10'd59) & ~(trunc_ln321_fu_8559_p1 == 10'd58) & ~(trunc_ln321_fu_8559_p1 == 10'd57) & ~(trunc_ln321_fu_8559_p1 == 10'd56) & ~(trunc_ln321_fu_8559_p1 == 10'd55) & ~(trunc_ln321_fu_8559_p1 == 10'd54) & ~(trunc_ln321_fu_8559_p1 == 10'd53) & ~(trunc_ln321_fu_8559_p1 == 10'd52) & ~(trunc_ln321_fu_8559_p1 == 10'd51) & ~(trunc_ln321_fu_8559_p1 == 10'd50) & ~(trunc_ln321_fu_8559_p1 == 10'd49) & ~(trunc_ln321_fu_8559_p1 == 10'd48) & ~(trunc_ln321_fu_8559_p1 == 10'd47) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd574) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd573) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd572) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd571) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd570) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd569) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd568) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd567) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd566) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd565) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd564) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd563) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd562) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd561) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd560) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd559) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd558) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd557) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd556) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd555) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd554) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd553) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd552) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd551) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd550) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd549) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd548) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd547) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd546) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd545) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd544) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd543) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd542) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd541) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd540) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd539) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd538) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd537) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd536) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd535) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd534) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd533) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd532) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd531) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd530) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd529) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd528) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd527) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd526) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd525) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd524) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd523) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd522) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd521) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd520) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd519) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd518) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd517) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd516) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd515) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd514) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd513) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd512) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd511) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd510) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd509) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd508) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd507) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd506) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd505) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd504) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd503) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd502) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd501) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd500) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd499) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd498) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd497) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd496) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd495) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd494) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd493) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd492) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd491) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd490) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd489) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd488) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd487) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd486) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd485) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd484) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd483) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd482) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd481) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd480) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd479) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd478) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd477) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd476) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd475) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd474) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd473) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd472) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd471) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd470) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd469) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd468) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd467) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd466) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd465) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd464) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd463) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd462) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd461) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd460) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd459) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd458) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd457) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd456) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd455) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd454) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd453) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd452) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd451) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd450) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd449) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd448) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd447) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd446) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd445) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd444) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd443) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd442) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd441) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd440) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd439) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd438) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd437) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd436) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd435) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd434) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd433) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd432) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd431) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd430) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd429) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd428) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd427) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd426) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd425) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd424) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd423) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd422) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd421) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd420) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd419) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd418) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd417) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd416) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd415) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd414) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd413) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd412) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd411) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd410) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd409) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd408) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd407) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd406) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd405) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd404) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd403) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd402) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd401) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd400) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd399) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd398) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd397) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd396) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd395) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd394) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd393) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd392) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd391) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd390) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd389) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd388) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd387) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd386) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd385) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd384) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd383) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd382) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd381) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd380) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd379) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd378) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd377) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd376) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd375) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd374) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd373) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd372) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd371) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd370) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd369) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd368) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd367) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd366) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd365) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd364) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd363) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd362) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd361) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd360) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd359) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd358) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd357) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd356) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd355) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd354) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd353) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd352) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd351) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd350) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd349) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd348) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd347) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd346) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd345) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd344) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd343) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd342) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd341) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd340) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd339) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd338) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd337) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd336) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd335) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd334) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd333) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd332) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd331) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd330) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd329) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd328) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd327) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd326) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd325) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd324) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd323) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd322) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd321) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd320) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd319) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd318) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd317) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd316) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd315) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd314) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd313) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd312) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd311) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd310) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd309) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd308) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd307) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd306) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd305) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd304) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd303) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd302) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd301) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd300) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd299) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd298) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd297) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd296) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd295) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd294) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd293) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd292) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd291) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd290) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd289) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd288) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd287) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd286) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd285) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd284) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd283) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd282) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd281) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd280) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd279) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd278) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd277) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd276) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd275) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd274) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd273) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd272) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd271) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd270) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd269) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd268) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd267) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd266) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd265) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd264) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd263) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd262) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd261) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd260) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd259) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd258) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd257) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd256) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd255) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd254) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd253) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd252) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd251) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd250) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd249) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd248) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd247) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd246) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd245) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd244) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd243) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd242) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd241) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd240) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd239) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd238) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd237) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd236) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd235) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd234) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd233) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd232) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd231) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd230) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd229) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd228) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd227) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd226) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd225) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd224) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd223) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd222) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd221) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd220) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd219) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd218) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd217) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd216) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd215) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd214) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd213) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd212) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd211) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd210) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd209) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd208) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd207) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd206) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd205) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd204) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd203) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd202) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd201) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd200) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd199) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd198) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd197) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd196) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd195) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd194) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd193) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd192) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd191) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd190) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd189) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd188) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd187) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd186) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd185) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd184) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd183) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd182) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd181) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd180) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd179) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd178) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd177) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd176) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd175) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd174) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd173) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd172) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd171) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd170) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd169) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd168) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd167) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd166) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd165) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd164) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd163) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd162) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd161) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd160) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd159) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd158) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd157) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd156) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd155) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd154) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd153) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd152) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd151) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd150) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd149) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd148) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd147) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd146) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd145) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd144) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd143) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd142) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd141) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd140) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd139) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd138) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd137) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd136) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd135) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd134) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd133) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd132) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd131) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd130) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd129) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd128) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd127) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd126) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd125) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd124) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd123) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd122) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd121) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd120) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd119) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd118) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd117) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd116) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd115) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd114) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd113) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd112) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd111) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd110) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd109) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd108) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd107) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd106) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd105) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd104) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd103) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd102) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd101) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd100) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd99) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd98) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd97) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd96) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd95) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd94) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd93) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd92) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd91) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd90) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd89) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd88) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd87) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd86) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd85) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd84) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd83) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd82) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd81) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd80) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd79) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd78) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd77) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd76) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd75) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd74) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd73) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd72) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd71) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd70) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd69) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd68) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd67) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd66) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd65) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd64) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd63) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd62) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd61) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd60) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd59) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd58) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd57) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd56) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd55) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd54) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd53) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd52) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd51) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd50) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd49) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd48) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((trunc_ln321_fu_8559_p1 == 10'd47) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_4476 <= in_V_V_TDATA;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_reg_pp0_iter1_act_m_val_V_reg_4476 <= ap_phi_reg_pp0_iter0_act_m_val_V_reg_4476;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_0_reg_4465 <= i_fu_5651_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_reg_4465 <= 16'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_17768 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        nf_assign_fu_3714 <= select_ln301_fu_11988_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        nf_assign_fu_3714 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_11612_p2 == 1'd0) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        sf_1_fu_1406 <= sf_fu_11606_p2;
    end else if ((((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_fu_11612_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        sf_1_fu_1406 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        accu_V_0_0_0_fu_1390 <= accu_0_0_V_fu_12053_p2;
        accu_V_0_1_0_fu_1394 <= accu_0_1_V_fu_12071_p2;
        accu_V_0_2_0_fu_1398 <= accu_0_2_V_fu_12089_p2;
        accu_V_0_3_0_fu_1402 <= accu_0_3_V_fu_12107_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln700_10_reg_17797 <= add_ln700_10_fu_11847_p2;
        add_ln700_14_reg_17807 <= add_ln700_14_fu_11907_p2;
        add_ln700_2_reg_17777 <= add_ln700_2_fu_11727_p2;
        add_ln700_6_reg_17787 <= add_ln700_6_fu_11787_p2;
        icmp_ln271_reg_17680_pp0_iter1_reg <= icmp_ln271_reg_17680;
        icmp_ln289_reg_17768_pp0_iter1_reg <= icmp_ln289_reg_17768;
        mul_ln1352_13_reg_17802 <= mul_ln1352_13_fu_11869_p2;
        mul_ln1352_1_reg_17772 <= mul_ln1352_1_fu_11661_p2;
        mul_ln1352_5_reg_17782 <= mul_ln1352_5_fu_11749_p2;
        mul_ln1352_9_reg_17792 <= mul_ln1352_9_fu_11809_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_5645_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln271_reg_17680 <= icmp_ln271_fu_11446_p2;
        icmp_ln289_reg_17768 <= icmp_ln289_fu_11612_p2;
        p_Result_1_0_1_reg_17693 <= {{weight_V_V_TDATA[7:4]}};
        p_Result_1_0_2_reg_17698 <= {{weight_V_V_TDATA[11:8]}};
        p_Result_1_0_3_reg_17703 <= {{weight_V_V_TDATA[15:12]}};
        p_Result_1_1_1_reg_17713 <= {{weight_V_V_TDATA[23:20]}};
        p_Result_1_1_2_reg_17718 <= {{weight_V_V_TDATA[27:24]}};
        p_Result_1_1_3_reg_17723 <= {{weight_V_V_TDATA[31:28]}};
        p_Result_1_1_reg_17708 <= {{weight_V_V_TDATA[19:16]}};
        p_Result_1_2_1_reg_17733 <= {{weight_V_V_TDATA[39:36]}};
        p_Result_1_2_2_reg_17738 <= {{weight_V_V_TDATA[43:40]}};
        p_Result_1_2_3_reg_17743 <= {{weight_V_V_TDATA[47:44]}};
        p_Result_1_2_reg_17728 <= {{weight_V_V_TDATA[35:32]}};
        p_Result_1_3_1_reg_17753 <= {{weight_V_V_TDATA[55:52]}};
        p_Result_1_3_2_reg_17758 <= {{weight_V_V_TDATA[59:56]}};
        p_Result_1_3_3_reg_17763 <= {{weight_V_V_TDATA[63:60]}};
        p_Result_1_3_reg_17748 <= {{weight_V_V_TDATA[51:48]}};
        trunc_ln647_reg_17688 <= trunc_ln647_fu_11452_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln289_reg_17768_pp0_iter2_reg <= icmp_ln289_reg_17768_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_17768_pp0_iter1_reg == 1'd1))) begin
        icmp_ln899_10_reg_18142 <= icmp_ln899_10_fu_12237_p2;
        icmp_ln899_11_reg_18147 <= icmp_ln899_11_fu_12247_p2;
        icmp_ln899_12_reg_18152 <= icmp_ln899_12_fu_12257_p2;
        icmp_ln899_13_reg_18157 <= icmp_ln899_13_fu_12267_p2;
        icmp_ln899_14_reg_18162 <= icmp_ln899_14_fu_12273_p2;
        icmp_ln899_15_reg_18167 <= icmp_ln899_15_fu_12279_p2;
        icmp_ln899_16_reg_18172 <= icmp_ln899_16_fu_12285_p2;
        icmp_ln899_17_reg_18177 <= icmp_ln899_17_fu_12291_p2;
        icmp_ln899_18_reg_18182 <= icmp_ln899_18_fu_12297_p2;
        icmp_ln899_19_reg_18187 <= icmp_ln899_19_fu_12303_p2;
        icmp_ln899_1_reg_18097 <= icmp_ln899_1_fu_12147_p2;
        icmp_ln899_20_reg_18192 <= icmp_ln899_20_fu_12309_p2;
        icmp_ln899_21_reg_18197 <= icmp_ln899_21_fu_12315_p2;
        icmp_ln899_22_reg_18202 <= icmp_ln899_22_fu_12321_p2;
        icmp_ln899_23_reg_18207 <= icmp_ln899_23_fu_12327_p2;
        icmp_ln899_24_reg_18212 <= icmp_ln899_24_fu_12333_p2;
        icmp_ln899_25_reg_18217 <= icmp_ln899_25_fu_12339_p2;
        icmp_ln899_26_reg_18222 <= icmp_ln899_26_fu_12345_p2;
        icmp_ln899_27_reg_18227 <= icmp_ln899_27_fu_12351_p2;
        icmp_ln899_28_reg_18232 <= icmp_ln899_28_fu_12361_p2;
        icmp_ln899_29_reg_18237 <= icmp_ln899_29_fu_12371_p2;
        icmp_ln899_2_reg_18102 <= icmp_ln899_2_fu_12157_p2;
        icmp_ln899_30_reg_18242 <= icmp_ln899_30_fu_12381_p2;
        icmp_ln899_31_reg_18247 <= icmp_ln899_31_fu_12391_p2;
        icmp_ln899_32_reg_18252 <= icmp_ln899_32_fu_12401_p2;
        icmp_ln899_33_reg_18257 <= icmp_ln899_33_fu_12411_p2;
        icmp_ln899_34_reg_18262 <= icmp_ln899_34_fu_12421_p2;
        icmp_ln899_35_reg_18267 <= icmp_ln899_35_fu_12431_p2;
        icmp_ln899_36_reg_18272 <= icmp_ln899_36_fu_12441_p2;
        icmp_ln899_37_reg_18277 <= icmp_ln899_37_fu_12451_p2;
        icmp_ln899_38_reg_18282 <= icmp_ln899_38_fu_12461_p2;
        icmp_ln899_39_reg_18287 <= icmp_ln899_39_fu_12471_p2;
        icmp_ln899_3_reg_18107 <= icmp_ln899_3_fu_12167_p2;
        icmp_ln899_40_reg_18292 <= icmp_ln899_40_fu_12481_p2;
        icmp_ln899_41_reg_18297 <= icmp_ln899_41_fu_12491_p2;
        icmp_ln899_42_reg_18302 <= icmp_ln899_42_fu_12497_p2;
        icmp_ln899_43_reg_18307 <= icmp_ln899_43_fu_12507_p2;
        icmp_ln899_44_reg_18312 <= icmp_ln899_44_fu_12517_p2;
        icmp_ln899_45_reg_18317 <= icmp_ln899_45_fu_12527_p2;
        icmp_ln899_46_reg_18322 <= icmp_ln899_46_fu_12537_p2;
        icmp_ln899_47_reg_18327 <= icmp_ln899_47_fu_12547_p2;
        icmp_ln899_48_reg_18332 <= icmp_ln899_48_fu_12557_p2;
        icmp_ln899_49_reg_18337 <= icmp_ln899_49_fu_12567_p2;
        icmp_ln899_4_reg_18112 <= icmp_ln899_4_fu_12177_p2;
        icmp_ln899_50_reg_18342 <= icmp_ln899_50_fu_12577_p2;
        icmp_ln899_51_reg_18347 <= icmp_ln899_51_fu_12587_p2;
        icmp_ln899_52_reg_18352 <= icmp_ln899_52_fu_12597_p2;
        icmp_ln899_53_reg_18357 <= icmp_ln899_53_fu_12607_p2;
        icmp_ln899_54_reg_18362 <= icmp_ln899_54_fu_12613_p2;
        icmp_ln899_55_reg_18367 <= icmp_ln899_55_fu_12619_p2;
        icmp_ln899_5_reg_18117 <= icmp_ln899_5_fu_12187_p2;
        icmp_ln899_6_reg_18122 <= icmp_ln899_6_fu_12197_p2;
        icmp_ln899_7_reg_18127 <= icmp_ln899_7_fu_12207_p2;
        icmp_ln899_8_reg_18132 <= icmp_ln899_8_fu_12217_p2;
        icmp_ln899_9_reg_18137 <= icmp_ln899_9_fu_12227_p2;
        icmp_ln899_reg_18092 <= icmp_ln899_fu_12137_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd99) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_100_fu_1806 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd100) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_101_fu_1810 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd101) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_102_fu_1814 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd102) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_103_fu_1818 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd103) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_104_fu_1822 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd104) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_105_fu_1826 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd105) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_106_fu_1830 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd106) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_107_fu_1834 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd107) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_108_fu_1838 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd108) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_109_fu_1842 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd9) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_10_fu_1446 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd109) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_110_fu_1846 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd110) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_111_fu_1850 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd111) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_112_fu_1854 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd112) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_113_fu_1858 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd113) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_114_fu_1862 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd114) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_115_fu_1866 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd115) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_116_fu_1870 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd116) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_117_fu_1874 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd117) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_118_fu_1878 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd118) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_119_fu_1882 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd10) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_11_fu_1450 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd119) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_120_fu_1886 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd120) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_121_fu_1890 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd121) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_122_fu_1894 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd122) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_123_fu_1898 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd123) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_124_fu_1902 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd124) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_125_fu_1906 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd125) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_126_fu_1910 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd126) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_127_fu_1914 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd127) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_128_fu_1918 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd128) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_129_fu_1922 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd11) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_12_fu_1454 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd129) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_130_fu_1926 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd130) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_131_fu_1930 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd131) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_132_fu_1934 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd132) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_133_fu_1938 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd133) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_134_fu_1942 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd134) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_135_fu_1946 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd135) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_136_fu_1950 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd136) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_137_fu_1954 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd137) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_138_fu_1958 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd138) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_139_fu_1962 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd12) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_13_fu_1458 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd139) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_140_fu_1966 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd140) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_141_fu_1970 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd141) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_142_fu_1974 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd142) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_143_fu_1978 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd143) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_144_fu_1982 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd144) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_145_fu_1986 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd145) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_146_fu_1990 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd146) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_147_fu_1994 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd147) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_148_fu_1998 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd148) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_149_fu_2002 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd13) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_14_fu_1462 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd149) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_150_fu_2006 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd150) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_151_fu_2010 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd151) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_152_fu_2014 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd152) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_153_fu_2018 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd153) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_154_fu_2022 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd154) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_155_fu_2026 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd155) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_156_fu_2030 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd156) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_157_fu_2034 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd157) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_158_fu_2038 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd158) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_159_fu_2042 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd14) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_15_fu_1466 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd159) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_160_fu_2046 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd160) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_161_fu_2050 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd161) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_162_fu_2054 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd162) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_163_fu_2058 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd163) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_164_fu_2062 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd164) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_165_fu_2066 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd165) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_166_fu_2070 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd166) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_167_fu_2074 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd167) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_168_fu_2078 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd168) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_169_fu_2082 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd15) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_16_fu_1470 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd169) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_170_fu_2086 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd170) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_171_fu_2090 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd171) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_172_fu_2094 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd172) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_173_fu_2098 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd173) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_174_fu_2102 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd174) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_175_fu_2106 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd175) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_176_fu_2110 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd176) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_177_fu_2114 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd177) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_178_fu_2118 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd178) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_179_fu_2122 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd16) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_17_fu_1474 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd179) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_180_fu_2126 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd180) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_181_fu_2130 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd181) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_182_fu_2134 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd182) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_183_fu_2138 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd183) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_184_fu_2142 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd184) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_185_fu_2146 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd185) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_186_fu_2150 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd186) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_187_fu_2154 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd187) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_188_fu_2158 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd188) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_189_fu_2162 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd17) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_18_fu_1478 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd189) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_190_fu_2166 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd190) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_191_fu_2170 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd191) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_192_fu_2174 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd192) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_193_fu_2178 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd193) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_194_fu_2182 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd194) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_195_fu_2186 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd195) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_196_fu_2190 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd196) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_197_fu_2194 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd197) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_198_fu_2198 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd198) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_199_fu_2202 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd18) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_19_fu_1482 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_1_fu_1414 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd199) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_200_fu_2206 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd200) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_201_fu_2210 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd201) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_202_fu_2214 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd202) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_203_fu_2218 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd203) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_204_fu_2222 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd204) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_205_fu_2226 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd205) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_206_fu_2230 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd206) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_207_fu_2234 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd207) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_208_fu_2238 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd208) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_209_fu_2242 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd19) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_20_fu_1486 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd209) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_210_fu_2246 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd210) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_211_fu_2250 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd211) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_212_fu_2254 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd212) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_213_fu_2258 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd213) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_214_fu_2262 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd214) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_215_fu_2266 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd215) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_216_fu_2270 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd216) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_217_fu_2274 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd217) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_218_fu_2278 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd218) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_219_fu_2282 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd20) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_21_fu_1490 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd219) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_220_fu_2286 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd220) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_221_fu_2290 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd221) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_222_fu_2294 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd222) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_223_fu_2298 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd223) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_224_fu_2302 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd224) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_225_fu_2306 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd225) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_226_fu_2310 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd226) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_227_fu_2314 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd227) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_228_fu_2318 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd228) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_229_fu_2322 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd21) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_22_fu_1494 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd229) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_230_fu_2326 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd230) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_231_fu_2330 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd231) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_232_fu_2334 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd232) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_233_fu_2338 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd233) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_234_fu_2342 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd234) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_235_fu_2346 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd235) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_236_fu_2350 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd236) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_237_fu_2354 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd237) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_238_fu_2358 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd238) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_239_fu_2362 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd22) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_23_fu_1498 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd239) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_240_fu_2366 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd240) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_241_fu_2370 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd241) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_242_fu_2374 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd242) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_243_fu_2378 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd243) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_244_fu_2382 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd244) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_245_fu_2386 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd245) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_246_fu_2390 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd246) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_247_fu_2394 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd247) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_248_fu_2398 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd248) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_249_fu_2402 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd23) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_24_fu_1502 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd249) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_250_fu_2406 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd250) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_251_fu_2410 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd251) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_252_fu_2414 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd252) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_253_fu_2418 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd253) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_254_fu_2422 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd254) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_255_fu_2426 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd255) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_256_fu_2430 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd256) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_257_fu_2434 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd257) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_258_fu_2438 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd258) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_259_fu_2442 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd24) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_25_fu_1506 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd259) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_260_fu_2446 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd260) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_261_fu_2450 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd261) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_262_fu_2454 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd262) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_263_fu_2458 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd263) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_264_fu_2462 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd264) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_265_fu_2466 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd265) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_266_fu_2470 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd266) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_267_fu_2474 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd267) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_268_fu_2478 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd268) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_269_fu_2482 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd25) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_26_fu_1510 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd269) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_270_fu_2486 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd270) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_271_fu_2490 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd271) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_272_fu_2494 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd272) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_273_fu_2498 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd273) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_274_fu_2502 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd274) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_275_fu_2506 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd275) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_276_fu_2510 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd276) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_277_fu_2514 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd277) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_278_fu_2518 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd278) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_279_fu_2522 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd26) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_27_fu_1514 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd279) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_280_fu_2526 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd280) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_281_fu_2530 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd281) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_282_fu_2534 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd282) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_283_fu_2538 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd283) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_284_fu_2542 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd284) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_285_fu_2546 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd285) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_286_fu_2550 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd286) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_287_fu_2554 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd287) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_288_fu_2558 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd288) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_289_fu_2562 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd27) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_28_fu_1518 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd289) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_290_fu_2566 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd290) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_291_fu_2570 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd291) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_292_fu_2574 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd292) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_293_fu_2578 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd293) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_294_fu_2582 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd294) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_295_fu_2586 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd295) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_296_fu_2590 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd296) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_297_fu_2594 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd297) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_298_fu_2598 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd298) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_299_fu_2602 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd28) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_29_fu_1522 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd2) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_2_fu_1418 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd299) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_300_fu_2606 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd300) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_301_fu_2610 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd301) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_302_fu_2614 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd302) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_303_fu_2618 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd303) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_304_fu_2622 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd304) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_305_fu_2626 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd305) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_306_fu_2630 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd306) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_307_fu_2634 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd307) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_308_fu_2638 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd308) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_309_fu_2642 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd29) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_30_fu_1526 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd309) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_310_fu_2646 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd310) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_311_fu_2650 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd311) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_312_fu_2654 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd312) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_313_fu_2658 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd313) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_314_fu_2662 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd314) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_315_fu_2666 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd315) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_316_fu_2670 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd316) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_317_fu_2674 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd317) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_318_fu_2678 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd318) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_319_fu_2682 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd30) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_31_fu_1530 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd319) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_320_fu_2686 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd320) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_321_fu_2690 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd321) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_322_fu_2694 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd322) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_323_fu_2698 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd323) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_324_fu_2702 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd324) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_325_fu_2706 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd325) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_326_fu_2710 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd326) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_327_fu_2714 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd327) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_328_fu_2718 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd328) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_329_fu_2722 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd31) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_32_fu_1534 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd329) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_330_fu_2726 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd330) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_331_fu_2730 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd331) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_332_fu_2734 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd332) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_333_fu_2738 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd333) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_334_fu_2742 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd334) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_335_fu_2746 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd335) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_336_fu_2750 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd336) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_337_fu_2754 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd337) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_338_fu_2758 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd338) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_339_fu_2762 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd32) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_33_fu_1538 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd339) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_340_fu_2766 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd340) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_341_fu_2770 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd341) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_342_fu_2774 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd342) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_343_fu_2778 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd343) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_344_fu_2782 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd344) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_345_fu_2786 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd345) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_346_fu_2790 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd346) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_347_fu_2794 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd347) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_348_fu_2798 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd348) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_349_fu_2802 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd33) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_34_fu_1542 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd349) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_350_fu_2806 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd350) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_351_fu_2810 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd351) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_352_fu_2814 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd352) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_353_fu_2818 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd353) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_354_fu_2822 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd354) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_355_fu_2826 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd355) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_356_fu_2830 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd356) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_357_fu_2834 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd357) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_358_fu_2838 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd358) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_359_fu_2842 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd34) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_35_fu_1546 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd359) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_360_fu_2846 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd360) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_361_fu_2850 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd361) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_362_fu_2854 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd362) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_363_fu_2858 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd363) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_364_fu_2862 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd364) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_365_fu_2866 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd365) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_366_fu_2870 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd366) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_367_fu_2874 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd367) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_368_fu_2878 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd368) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_369_fu_2882 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd35) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_36_fu_1550 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd369) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_370_fu_2886 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd370) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_371_fu_2890 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd371) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_372_fu_2894 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd372) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_373_fu_2898 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd373) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_374_fu_2902 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd374) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_375_fu_2906 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd375) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_376_fu_2910 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd376) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_377_fu_2914 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd377) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_378_fu_2918 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd378) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_379_fu_2922 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd36) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_37_fu_1554 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd379) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_380_fu_2926 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd380) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_381_fu_2930 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd381) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_382_fu_2934 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd382) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_383_fu_2938 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd383) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_384_fu_2942 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd384) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_385_fu_2946 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd385) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_386_fu_2950 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd386) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_387_fu_2954 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd387) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_388_fu_2958 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd388) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_389_fu_2962 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd37) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_38_fu_1558 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd389) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_390_fu_2966 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd390) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_391_fu_2970 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd391) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_392_fu_2974 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd392) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_393_fu_2978 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd393) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_394_fu_2982 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd394) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_395_fu_2986 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd395) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_396_fu_2990 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd396) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_397_fu_2994 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd397) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_398_fu_2998 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd398) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_399_fu_3002 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd38) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_39_fu_1562 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd399) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_400_fu_3006 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd400) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_401_fu_3010 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd401) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_402_fu_3014 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd402) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_403_fu_3018 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd403) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_404_fu_3022 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd404) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_405_fu_3026 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd405) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_406_fu_3030 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd406) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_407_fu_3034 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd407) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_408_fu_3038 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd408) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_409_fu_3042 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd39) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_40_fu_1566 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd409) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_410_fu_3046 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd410) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_411_fu_3050 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd411) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_412_fu_3054 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd412) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_413_fu_3058 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd413) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_414_fu_3062 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd414) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_415_fu_3066 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd415) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_416_fu_3070 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd416) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_417_fu_3074 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd417) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_418_fu_3078 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd418) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_419_fu_3082 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd40) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_41_fu_1570 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd419) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_420_fu_3086 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd420) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_421_fu_3090 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd421) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_422_fu_3094 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd422) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_423_fu_3098 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd423) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_424_fu_3102 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd424) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_425_fu_3106 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd425) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_426_fu_3110 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd426) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_427_fu_3114 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd427) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_428_fu_3118 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd428) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_429_fu_3122 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd41) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_42_fu_1574 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd429) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_430_fu_3126 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd430) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_431_fu_3130 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd431) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_432_fu_3134 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd432) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_433_fu_3138 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd433) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_434_fu_3142 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd434) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_435_fu_3146 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd435) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_436_fu_3150 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd436) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_437_fu_3154 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd437) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_438_fu_3158 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd438) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_439_fu_3162 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd42) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_43_fu_1578 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd439) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_440_fu_3166 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd440) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_441_fu_3170 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd441) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_442_fu_3174 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd442) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_443_fu_3178 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd443) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_444_fu_3182 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd444) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_445_fu_3186 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd445) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_446_fu_3190 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd446) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_447_fu_3194 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd447) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_448_fu_3198 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd448) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_449_fu_3202 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd43) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_44_fu_1582 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd449) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_450_fu_3206 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd450) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_451_fu_3210 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd451) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_452_fu_3214 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd452) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_453_fu_3218 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd453) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_454_fu_3222 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd454) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_455_fu_3226 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd455) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_456_fu_3230 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd456) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_457_fu_3234 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd457) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_458_fu_3238 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd458) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_459_fu_3242 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd44) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_45_fu_1586 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd459) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_460_fu_3246 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd460) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_461_fu_3250 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd461) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_462_fu_3254 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd462) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_463_fu_3258 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd463) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_464_fu_3262 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd464) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_465_fu_3266 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd465) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_466_fu_3270 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd466) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_467_fu_3274 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd467) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_468_fu_3278 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd468) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_469_fu_3282 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd45) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_46_fu_1590 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd469) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_470_fu_3286 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd470) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_471_fu_3290 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd471) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_472_fu_3294 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd472) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_473_fu_3298 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd473) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_474_fu_3302 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd474) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_475_fu_3306 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd475) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_476_fu_3310 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd476) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_477_fu_3314 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd477) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_478_fu_3318 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd478) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_479_fu_3322 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd46) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_47_fu_1594 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd479) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_480_fu_3326 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd480) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_481_fu_3330 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd481) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_482_fu_3334 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd482) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_483_fu_3338 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd483) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_484_fu_3342 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd484) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_485_fu_3346 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd485) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_486_fu_3350 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd486) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_487_fu_3354 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd487) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_488_fu_3358 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd488) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_489_fu_3362 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd47) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_48_fu_1598 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd489) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_490_fu_3366 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd490) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_491_fu_3370 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd491) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_492_fu_3374 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd492) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_493_fu_3378 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd493) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_494_fu_3382 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd494) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_495_fu_3386 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd495) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_496_fu_3390 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd496) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_497_fu_3394 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd497) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_498_fu_3398 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd498) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_499_fu_3402 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd48) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_49_fu_1602 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd3) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_4_fu_1422 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd499) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_500_fu_3406 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd500) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_501_fu_3410 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd501) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_502_fu_3414 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd502) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_503_fu_3418 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd503) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_504_fu_3422 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd504) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_505_fu_3426 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd505) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_506_fu_3430 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd506) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_507_fu_3434 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd507) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_508_fu_3438 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd508) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_509_fu_3442 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd49) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_50_fu_1606 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd509) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_510_fu_3446 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd510) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_511_fu_3450 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd511) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_512_fu_3454 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd512) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_513_fu_3458 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd513) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_514_fu_3462 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd514) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_515_fu_3466 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd515) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_516_fu_3470 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd516) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_517_fu_3474 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd517) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_518_fu_3478 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd518) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_519_fu_3482 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd50) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_51_fu_1610 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd519) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_520_fu_3486 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd520) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_521_fu_3490 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd521) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_522_fu_3494 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd522) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_523_fu_3498 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd523) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_524_fu_3502 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd524) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_525_fu_3506 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd525) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_526_fu_3510 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd526) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_527_fu_3514 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd527) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_528_fu_3518 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd528) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_529_fu_3522 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd51) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_52_fu_1614 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd529) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_530_fu_3526 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd530) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_531_fu_3530 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd531) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_532_fu_3534 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd532) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_533_fu_3538 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd533) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_534_fu_3542 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd534) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_535_fu_3546 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd535) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_536_fu_3550 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd536) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_537_fu_3554 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd537) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_538_fu_3558 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd538) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_539_fu_3562 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd52) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_53_fu_1618 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd539) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_540_fu_3566 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd540) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_541_fu_3570 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd541) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_542_fu_3574 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd542) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_543_fu_3578 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd543) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_544_fu_3582 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd544) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_545_fu_3586 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd545) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_546_fu_3590 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd546) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_547_fu_3594 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd547) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_548_fu_3598 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd548) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_549_fu_3602 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd53) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_54_fu_1622 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd549) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_550_fu_3606 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd550) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_551_fu_3610 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd551) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_552_fu_3614 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd552) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_553_fu_3618 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd553) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_554_fu_3622 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd554) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_555_fu_3626 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd555) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_556_fu_3630 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd556) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_557_fu_3634 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd557) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_558_fu_3638 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd558) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_559_fu_3642 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd54) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_55_fu_1626 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd559) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_560_fu_3646 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd560) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_561_fu_3650 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd561) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_562_fu_3654 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd562) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_563_fu_3658 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd563) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_564_fu_3662 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd564) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_565_fu_3666 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd565) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_566_fu_3670 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd566) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_567_fu_3674 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd567) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_568_fu_3678 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd568) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_569_fu_3682 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd55) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_56_fu_1630 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd569) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_570_fu_3686 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd570) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_571_fu_3690 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd571) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_572_fu_3694 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd572) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_573_fu_3698 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd573) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_574_fu_3702 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd574) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_575_fu_3706 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if ((~(trunc_ln321_fu_8559_p1 == 10'd46) & ~(trunc_ln321_fu_8559_p1 == 10'd45) & ~(trunc_ln321_fu_8559_p1 == 10'd44) & ~(trunc_ln321_fu_8559_p1 == 10'd43) & ~(trunc_ln321_fu_8559_p1 == 10'd42) & ~(trunc_ln321_fu_8559_p1 == 10'd41) & ~(trunc_ln321_fu_8559_p1 == 10'd40) & ~(trunc_ln321_fu_8559_p1 == 10'd39) & ~(trunc_ln321_fu_8559_p1 == 10'd38) & ~(trunc_ln321_fu_8559_p1 == 10'd37) & ~(trunc_ln321_fu_8559_p1 == 10'd36) & ~(trunc_ln321_fu_8559_p1 == 10'd35) & ~(trunc_ln321_fu_8559_p1 == 10'd34) & ~(trunc_ln321_fu_8559_p1 == 10'd33) & ~(trunc_ln321_fu_8559_p1 == 10'd32) & ~(trunc_ln321_fu_8559_p1 == 10'd31) & ~(trunc_ln321_fu_8559_p1 == 10'd30) & ~(trunc_ln321_fu_8559_p1 == 10'd29) & ~(trunc_ln321_fu_8559_p1 == 10'd28) & ~(trunc_ln321_fu_8559_p1 == 10'd27) & ~(trunc_ln321_fu_8559_p1 == 10'd26) & ~(trunc_ln321_fu_8559_p1 == 10'd25) & ~(trunc_ln321_fu_8559_p1 == 10'd24) & ~(trunc_ln321_fu_8559_p1 == 10'd23) & ~(trunc_ln321_fu_8559_p1 == 10'd22) & ~(trunc_ln321_fu_8559_p1 == 10'd21) & ~(trunc_ln321_fu_8559_p1 == 10'd20) & ~(trunc_ln321_fu_8559_p1 == 10'd19) & ~(trunc_ln321_fu_8559_p1 == 10'd18) & ~(trunc_ln321_fu_8559_p1 == 10'd17) & ~(trunc_ln321_fu_8559_p1 == 10'd16) & ~(trunc_ln321_fu_8559_p1 == 10'd15) & ~(trunc_ln321_fu_8559_p1 == 10'd14) & ~(trunc_ln321_fu_8559_p1 == 10'd13) & ~(trunc_ln321_fu_8559_p1 == 10'd12) & ~(trunc_ln321_fu_8559_p1 == 10'd11) & ~(trunc_ln321_fu_8559_p1 == 10'd10) & ~(trunc_ln321_fu_8559_p1 == 10'd9) & ~(trunc_ln321_fu_8559_p1 == 10'd8) & ~(trunc_ln321_fu_8559_p1 == 10'd7) & ~(trunc_ln321_fu_8559_p1 == 10'd6) & ~(trunc_ln321_fu_8559_p1 == 10'd5) & ~(trunc_ln321_fu_8559_p1 == 10'd4) & ~(trunc_ln321_fu_8559_p1 == 10'd3) & ~(trunc_ln321_fu_8559_p1 == 10'd2) & ~(trunc_ln321_fu_8559_p1 == 10'd1) & ~(trunc_ln321_fu_8559_p1 == 10'd0) & ~(trunc_ln321_fu_8559_p1 == 10'd574) & ~(trunc_ln321_fu_8559_p1 == 10'd573) & ~(trunc_ln321_fu_8559_p1 == 10'd572) & ~(trunc_ln321_fu_8559_p1 == 10'd571) & ~(trunc_ln321_fu_8559_p1 == 10'd570) & ~(trunc_ln321_fu_8559_p1 == 10'd569) & ~(trunc_ln321_fu_8559_p1 == 10'd568) & ~(trunc_ln321_fu_8559_p1 == 10'd567) & ~(trunc_ln321_fu_8559_p1 == 10'd566) & ~(trunc_ln321_fu_8559_p1 == 10'd565) & ~(trunc_ln321_fu_8559_p1 == 10'd564) & ~(trunc_ln321_fu_8559_p1 == 10'd563) & ~(trunc_ln321_fu_8559_p1 == 10'd562) & ~(trunc_ln321_fu_8559_p1 == 10'd561) & ~(trunc_ln321_fu_8559_p1 == 10'd560) & ~(trunc_ln321_fu_8559_p1 == 10'd559) & ~(trunc_ln321_fu_8559_p1 == 10'd558) & ~(trunc_ln321_fu_8559_p1 == 10'd557) & ~(trunc_ln321_fu_8559_p1 == 10'd556) & ~(trunc_ln321_fu_8559_p1 == 10'd555) & ~(trunc_ln321_fu_8559_p1 == 10'd554) & ~(trunc_ln321_fu_8559_p1 == 10'd553) & ~(trunc_ln321_fu_8559_p1 == 10'd552) & ~(trunc_ln321_fu_8559_p1 == 10'd551) & ~(trunc_ln321_fu_8559_p1 == 10'd550) & ~(trunc_ln321_fu_8559_p1 == 10'd549) & ~(trunc_ln321_fu_8559_p1 == 10'd548) & ~(trunc_ln321_fu_8559_p1 == 10'd547) & ~(trunc_ln321_fu_8559_p1 == 10'd546) & ~(trunc_ln321_fu_8559_p1 == 10'd545) & ~(trunc_ln321_fu_8559_p1 == 10'd544) & ~(trunc_ln321_fu_8559_p1 == 10'd543) & ~(trunc_ln321_fu_8559_p1 == 10'd542) & ~(trunc_ln321_fu_8559_p1 == 10'd541) & ~(trunc_ln321_fu_8559_p1 == 10'd540) & ~(trunc_ln321_fu_8559_p1 == 10'd539) & ~(trunc_ln321_fu_8559_p1 == 10'd538) & ~(trunc_ln321_fu_8559_p1 == 10'd537) & ~(trunc_ln321_fu_8559_p1 == 10'd536) & ~(trunc_ln321_fu_8559_p1 == 10'd535) & ~(trunc_ln321_fu_8559_p1 == 10'd534) & ~(trunc_ln321_fu_8559_p1 == 10'd533) & ~(trunc_ln321_fu_8559_p1 == 10'd532) & ~(trunc_ln321_fu_8559_p1 == 10'd531) & ~(trunc_ln321_fu_8559_p1 == 10'd530) & ~(trunc_ln321_fu_8559_p1 == 10'd529) & ~(trunc_ln321_fu_8559_p1 == 10'd528) & ~(trunc_ln321_fu_8559_p1 == 10'd527) & ~(trunc_ln321_fu_8559_p1 == 10'd526) & ~(trunc_ln321_fu_8559_p1 == 10'd525) & ~(trunc_ln321_fu_8559_p1 == 10'd524) & ~(trunc_ln321_fu_8559_p1 == 10'd523) & ~(trunc_ln321_fu_8559_p1 == 10'd522) & ~(trunc_ln321_fu_8559_p1 == 10'd521) & ~(trunc_ln321_fu_8559_p1 == 10'd520) & ~(trunc_ln321_fu_8559_p1 == 10'd519) & ~(trunc_ln321_fu_8559_p1 == 10'd518) & ~(trunc_ln321_fu_8559_p1 == 10'd517) & ~(trunc_ln321_fu_8559_p1 == 10'd516) & ~(trunc_ln321_fu_8559_p1 == 10'd515) & ~(trunc_ln321_fu_8559_p1 == 10'd514) & ~(trunc_ln321_fu_8559_p1 == 10'd513) & ~(trunc_ln321_fu_8559_p1 == 10'd512) & ~(trunc_ln321_fu_8559_p1 == 10'd511) & ~(trunc_ln321_fu_8559_p1 == 10'd510) & ~(trunc_ln321_fu_8559_p1 == 10'd509) & ~(trunc_ln321_fu_8559_p1 == 10'd508) & ~(trunc_ln321_fu_8559_p1 == 10'd507) & ~(trunc_ln321_fu_8559_p1 == 10'd506) & ~(trunc_ln321_fu_8559_p1 == 10'd505) & ~(trunc_ln321_fu_8559_p1 == 10'd504) & ~(trunc_ln321_fu_8559_p1 == 10'd503) & ~(trunc_ln321_fu_8559_p1 == 10'd502) & ~(trunc_ln321_fu_8559_p1 == 10'd501) & ~(trunc_ln321_fu_8559_p1 == 10'd500) & ~(trunc_ln321_fu_8559_p1 == 10'd499) & ~(trunc_ln321_fu_8559_p1 == 10'd498) & ~(trunc_ln321_fu_8559_p1 == 10'd497) & ~(trunc_ln321_fu_8559_p1 == 10'd496) & ~(trunc_ln321_fu_8559_p1 == 10'd495) & ~(trunc_ln321_fu_8559_p1 == 10'd494) & ~(trunc_ln321_fu_8559_p1 == 10'd493) & ~(trunc_ln321_fu_8559_p1 == 10'd492) & ~(trunc_ln321_fu_8559_p1 == 10'd491) & ~(trunc_ln321_fu_8559_p1 == 10'd490) & ~(trunc_ln321_fu_8559_p1 == 10'd489) & ~(trunc_ln321_fu_8559_p1 == 10'd488) & ~(trunc_ln321_fu_8559_p1 == 10'd487) & ~(trunc_ln321_fu_8559_p1 == 10'd486) & ~(trunc_ln321_fu_8559_p1 == 10'd485) & ~(trunc_ln321_fu_8559_p1 == 10'd484) & ~(trunc_ln321_fu_8559_p1 == 10'd483) & ~(trunc_ln321_fu_8559_p1 == 10'd482) & ~(trunc_ln321_fu_8559_p1 == 10'd481) & ~(trunc_ln321_fu_8559_p1 == 10'd480) & ~(trunc_ln321_fu_8559_p1 == 10'd479) & ~(trunc_ln321_fu_8559_p1 == 10'd478) & ~(trunc_ln321_fu_8559_p1 == 10'd477) & ~(trunc_ln321_fu_8559_p1 == 10'd476) & ~(trunc_ln321_fu_8559_p1 == 10'd475) & ~(trunc_ln321_fu_8559_p1 == 10'd474) & ~(trunc_ln321_fu_8559_p1 == 10'd473) & ~(trunc_ln321_fu_8559_p1 == 10'd472) & ~(trunc_ln321_fu_8559_p1 == 10'd471) & ~(trunc_ln321_fu_8559_p1 == 10'd470) & ~(trunc_ln321_fu_8559_p1 == 10'd469) & ~(trunc_ln321_fu_8559_p1 == 10'd468) & ~(trunc_ln321_fu_8559_p1 == 10'd467) & ~(trunc_ln321_fu_8559_p1 == 10'd466) & ~(trunc_ln321_fu_8559_p1 == 10'd465) & ~(trunc_ln321_fu_8559_p1 == 10'd464) & ~(trunc_ln321_fu_8559_p1 == 10'd463) & ~(trunc_ln321_fu_8559_p1 == 10'd462) & ~(trunc_ln321_fu_8559_p1 == 10'd461) & ~(trunc_ln321_fu_8559_p1 == 10'd460) & ~(trunc_ln321_fu_8559_p1 == 10'd459) & ~(trunc_ln321_fu_8559_p1 == 10'd458) & ~(trunc_ln321_fu_8559_p1 == 10'd457) & ~(trunc_ln321_fu_8559_p1 == 10'd456) & ~(trunc_ln321_fu_8559_p1 == 10'd455) & ~(trunc_ln321_fu_8559_p1 == 10'd454) & ~(trunc_ln321_fu_8559_p1 == 10'd453) & ~(trunc_ln321_fu_8559_p1 == 10'd452) & ~(trunc_ln321_fu_8559_p1 == 10'd451) & ~(trunc_ln321_fu_8559_p1 == 10'd450) & ~(trunc_ln321_fu_8559_p1 == 10'd449) & ~(trunc_ln321_fu_8559_p1 == 10'd448) & ~(trunc_ln321_fu_8559_p1 == 10'd447) & ~(trunc_ln321_fu_8559_p1 == 10'd446) & ~(trunc_ln321_fu_8559_p1 == 10'd445) & ~(trunc_ln321_fu_8559_p1 == 10'd444) & ~(trunc_ln321_fu_8559_p1 == 10'd443) & ~(trunc_ln321_fu_8559_p1 == 10'd442) & ~(trunc_ln321_fu_8559_p1 == 10'd441) & ~(trunc_ln321_fu_8559_p1 == 10'd440) & ~(trunc_ln321_fu_8559_p1 == 10'd439) & ~(trunc_ln321_fu_8559_p1 == 10'd438) & ~(trunc_ln321_fu_8559_p1 == 10'd437) & ~(trunc_ln321_fu_8559_p1 == 10'd436) & ~(trunc_ln321_fu_8559_p1 == 10'd435) & ~(trunc_ln321_fu_8559_p1 == 10'd434) & ~(trunc_ln321_fu_8559_p1 == 10'd433) & ~(trunc_ln321_fu_8559_p1 == 10'd432) & ~(trunc_ln321_fu_8559_p1 == 10'd431) & ~(trunc_ln321_fu_8559_p1 == 10'd430) & ~(trunc_ln321_fu_8559_p1 == 10'd429) & ~(trunc_ln321_fu_8559_p1 == 10'd428) & ~(trunc_ln321_fu_8559_p1 == 10'd427) & ~(trunc_ln321_fu_8559_p1 == 10'd426) & ~(trunc_ln321_fu_8559_p1 == 10'd425) & ~(trunc_ln321_fu_8559_p1 == 10'd424) & ~(trunc_ln321_fu_8559_p1 == 10'd423) & ~(trunc_ln321_fu_8559_p1 == 10'd422) & ~(trunc_ln321_fu_8559_p1 == 10'd421) & ~(trunc_ln321_fu_8559_p1 == 10'd420) & ~(trunc_ln321_fu_8559_p1 == 10'd419) & ~(trunc_ln321_fu_8559_p1 == 10'd418) & ~(trunc_ln321_fu_8559_p1 == 10'd417) & ~(trunc_ln321_fu_8559_p1 == 10'd416) & ~(trunc_ln321_fu_8559_p1 == 10'd415) & ~(trunc_ln321_fu_8559_p1 == 10'd414) & ~(trunc_ln321_fu_8559_p1 == 10'd413) & ~(trunc_ln321_fu_8559_p1 == 10'd412) & ~(trunc_ln321_fu_8559_p1 == 10'd411) & ~(trunc_ln321_fu_8559_p1 == 10'd410) & ~(trunc_ln321_fu_8559_p1 == 10'd409) & ~(trunc_ln321_fu_8559_p1 == 10'd408) & ~(trunc_ln321_fu_8559_p1 == 10'd407) & ~(trunc_ln321_fu_8559_p1 == 10'd406) & ~(trunc_ln321_fu_8559_p1 == 10'd405) & ~(trunc_ln321_fu_8559_p1 == 10'd404) & ~(trunc_ln321_fu_8559_p1 == 10'd403) & ~(trunc_ln321_fu_8559_p1 == 10'd402) & ~(trunc_ln321_fu_8559_p1 == 10'd401) & ~(trunc_ln321_fu_8559_p1 == 10'd400) & ~(trunc_ln321_fu_8559_p1 == 10'd399) & ~(trunc_ln321_fu_8559_p1 == 10'd398) & ~(trunc_ln321_fu_8559_p1 == 10'd397) & ~(trunc_ln321_fu_8559_p1 == 10'd396) & ~(trunc_ln321_fu_8559_p1 == 10'd395) & ~(trunc_ln321_fu_8559_p1 == 10'd394) & ~(trunc_ln321_fu_8559_p1 == 10'd393) & ~(trunc_ln321_fu_8559_p1 == 10'd392) & ~(trunc_ln321_fu_8559_p1 == 10'd391) & ~(trunc_ln321_fu_8559_p1 == 10'd390) & ~(trunc_ln321_fu_8559_p1 == 10'd389) & ~(trunc_ln321_fu_8559_p1 == 10'd388) & ~(trunc_ln321_fu_8559_p1 == 10'd387) & ~(trunc_ln321_fu_8559_p1 == 10'd386) & ~(trunc_ln321_fu_8559_p1 == 10'd385) & ~(trunc_ln321_fu_8559_p1 == 10'd384) & ~(trunc_ln321_fu_8559_p1 == 10'd383) & ~(trunc_ln321_fu_8559_p1 == 10'd382) & ~(trunc_ln321_fu_8559_p1 == 10'd381) & ~(trunc_ln321_fu_8559_p1 == 10'd380) & ~(trunc_ln321_fu_8559_p1 == 10'd379) & ~(trunc_ln321_fu_8559_p1 == 10'd378) & ~(trunc_ln321_fu_8559_p1 == 10'd377) & ~(trunc_ln321_fu_8559_p1 == 10'd376) & ~(trunc_ln321_fu_8559_p1 == 10'd375) & ~(trunc_ln321_fu_8559_p1 == 10'd374) & ~(trunc_ln321_fu_8559_p1 == 10'd373) & ~(trunc_ln321_fu_8559_p1 == 10'd372) & ~(trunc_ln321_fu_8559_p1 == 10'd371) & ~(trunc_ln321_fu_8559_p1 == 10'd370) & ~(trunc_ln321_fu_8559_p1 == 10'd369) & ~(trunc_ln321_fu_8559_p1 == 10'd368) & ~(trunc_ln321_fu_8559_p1 == 10'd367) & ~(trunc_ln321_fu_8559_p1 == 10'd366) & ~(trunc_ln321_fu_8559_p1 == 10'd365) & ~(trunc_ln321_fu_8559_p1 == 10'd364) & ~(trunc_ln321_fu_8559_p1 == 10'd363) & ~(trunc_ln321_fu_8559_p1 == 10'd362) & ~(trunc_ln321_fu_8559_p1 == 10'd361) & ~(trunc_ln321_fu_8559_p1 == 10'd360) & ~(trunc_ln321_fu_8559_p1 == 10'd359) & ~(trunc_ln321_fu_8559_p1 == 10'd358) & ~(trunc_ln321_fu_8559_p1 == 10'd357) & ~(trunc_ln321_fu_8559_p1 == 10'd356) & ~(trunc_ln321_fu_8559_p1 == 10'd355) & ~(trunc_ln321_fu_8559_p1 == 10'd354) & ~(trunc_ln321_fu_8559_p1 == 10'd353) & ~(trunc_ln321_fu_8559_p1 == 10'd352) & ~(trunc_ln321_fu_8559_p1 == 10'd351) & ~(trunc_ln321_fu_8559_p1 == 10'd350) & ~(trunc_ln321_fu_8559_p1 == 10'd349) & ~(trunc_ln321_fu_8559_p1 == 10'd348) & ~(trunc_ln321_fu_8559_p1 == 10'd347) & ~(trunc_ln321_fu_8559_p1 == 10'd346) & ~(trunc_ln321_fu_8559_p1 == 10'd345) & ~(trunc_ln321_fu_8559_p1 == 10'd344) & ~(trunc_ln321_fu_8559_p1 == 10'd343) & ~(trunc_ln321_fu_8559_p1 == 10'd342) & ~(trunc_ln321_fu_8559_p1 == 10'd341) & ~(trunc_ln321_fu_8559_p1 == 10'd340) & ~(trunc_ln321_fu_8559_p1 == 10'd339) & ~(trunc_ln321_fu_8559_p1 == 10'd338) & ~(trunc_ln321_fu_8559_p1 == 10'd337) & ~(trunc_ln321_fu_8559_p1 == 10'd336) & ~(trunc_ln321_fu_8559_p1 == 10'd335) & ~(trunc_ln321_fu_8559_p1 == 10'd334) & ~(trunc_ln321_fu_8559_p1 == 10'd333) & ~(trunc_ln321_fu_8559_p1 == 10'd332) & ~(trunc_ln321_fu_8559_p1 == 10'd331) & ~(trunc_ln321_fu_8559_p1 == 10'd330) & ~(trunc_ln321_fu_8559_p1 == 10'd329) & ~(trunc_ln321_fu_8559_p1 == 10'd328) & ~(trunc_ln321_fu_8559_p1 == 10'd327) & ~(trunc_ln321_fu_8559_p1 == 10'd326) & ~(trunc_ln321_fu_8559_p1 == 10'd325) & ~(trunc_ln321_fu_8559_p1 == 10'd324) & ~(trunc_ln321_fu_8559_p1 == 10'd323) & ~(trunc_ln321_fu_8559_p1 == 10'd322) & ~(trunc_ln321_fu_8559_p1 == 10'd321) & ~(trunc_ln321_fu_8559_p1 == 10'd320) & ~(trunc_ln321_fu_8559_p1 == 10'd319) & ~(trunc_ln321_fu_8559_p1 == 10'd318) & ~(trunc_ln321_fu_8559_p1 == 10'd317) & ~(trunc_ln321_fu_8559_p1 == 10'd316) & ~(trunc_ln321_fu_8559_p1 == 10'd315) & ~(trunc_ln321_fu_8559_p1 == 10'd314) & ~(trunc_ln321_fu_8559_p1 == 10'd313) & ~(trunc_ln321_fu_8559_p1 == 10'd312) & ~(trunc_ln321_fu_8559_p1 == 10'd311) & ~(trunc_ln321_fu_8559_p1 == 10'd310) & ~(trunc_ln321_fu_8559_p1 == 10'd309) & ~(trunc_ln321_fu_8559_p1 == 10'd308) & ~(trunc_ln321_fu_8559_p1 == 10'd307) & ~(trunc_ln321_fu_8559_p1 == 10'd306) & ~(trunc_ln321_fu_8559_p1 == 10'd305) & ~(trunc_ln321_fu_8559_p1 == 10'd304) & ~(trunc_ln321_fu_8559_p1 == 10'd303) & ~(trunc_ln321_fu_8559_p1 == 10'd302) & ~(trunc_ln321_fu_8559_p1 == 10'd301) & ~(trunc_ln321_fu_8559_p1 == 10'd300) & ~(trunc_ln321_fu_8559_p1 == 10'd299) & ~(trunc_ln321_fu_8559_p1 == 10'd298) & ~(trunc_ln321_fu_8559_p1 == 10'd297) & ~(trunc_ln321_fu_8559_p1 == 10'd296) & ~(trunc_ln321_fu_8559_p1 == 10'd295) & ~(trunc_ln321_fu_8559_p1 == 10'd294) & ~(trunc_ln321_fu_8559_p1 == 10'd293) & ~(trunc_ln321_fu_8559_p1 == 10'd292) & ~(trunc_ln321_fu_8559_p1 == 10'd291) & ~(trunc_ln321_fu_8559_p1 == 10'd290) & ~(trunc_ln321_fu_8559_p1 == 10'd289) & ~(trunc_ln321_fu_8559_p1 == 10'd288) & ~(trunc_ln321_fu_8559_p1 == 10'd287) & ~(trunc_ln321_fu_8559_p1 == 10'd286) & ~(trunc_ln321_fu_8559_p1 == 10'd285) & ~(trunc_ln321_fu_8559_p1 == 10'd284) & ~(trunc_ln321_fu_8559_p1 == 10'd283) & ~(trunc_ln321_fu_8559_p1 == 10'd282) & ~(trunc_ln321_fu_8559_p1 == 10'd281) & ~(trunc_ln321_fu_8559_p1 == 10'd280) & ~(trunc_ln321_fu_8559_p1 == 10'd279) & ~(trunc_ln321_fu_8559_p1 == 10'd278) & ~(trunc_ln321_fu_8559_p1 == 10'd277) & ~(trunc_ln321_fu_8559_p1 == 10'd276) & ~(trunc_ln321_fu_8559_p1 == 10'd275) & ~(trunc_ln321_fu_8559_p1 == 10'd274) & ~(trunc_ln321_fu_8559_p1 == 10'd273) & ~(trunc_ln321_fu_8559_p1 == 10'd272) & ~(trunc_ln321_fu_8559_p1 == 10'd271) & ~(trunc_ln321_fu_8559_p1 == 10'd270) & ~(trunc_ln321_fu_8559_p1 == 10'd269) & ~(trunc_ln321_fu_8559_p1 == 10'd268) & ~(trunc_ln321_fu_8559_p1 == 10'd267) & ~(trunc_ln321_fu_8559_p1 == 10'd266) & ~(trunc_ln321_fu_8559_p1 == 10'd265) & ~(trunc_ln321_fu_8559_p1 == 10'd264) & ~(trunc_ln321_fu_8559_p1 == 10'd263) & ~(trunc_ln321_fu_8559_p1 == 10'd262) & ~(trunc_ln321_fu_8559_p1 == 10'd261) & ~(trunc_ln321_fu_8559_p1 == 10'd260) & ~(trunc_ln321_fu_8559_p1 == 10'd259) & ~(trunc_ln321_fu_8559_p1 == 10'd258) & ~(trunc_ln321_fu_8559_p1 == 10'd257) & ~(trunc_ln321_fu_8559_p1 == 10'd256) & ~(trunc_ln321_fu_8559_p1 == 10'd255) & ~(trunc_ln321_fu_8559_p1 == 10'd254) & ~(trunc_ln321_fu_8559_p1 == 10'd253) & ~(trunc_ln321_fu_8559_p1 == 10'd252) & ~(trunc_ln321_fu_8559_p1 == 10'd251) & ~(trunc_ln321_fu_8559_p1 == 10'd250) & ~(trunc_ln321_fu_8559_p1 == 10'd249) & ~(trunc_ln321_fu_8559_p1 == 10'd248) & ~(trunc_ln321_fu_8559_p1 == 10'd247) & ~(trunc_ln321_fu_8559_p1 == 10'd246) & ~(trunc_ln321_fu_8559_p1 == 10'd245) & ~(trunc_ln321_fu_8559_p1 == 10'd244) & ~(trunc_ln321_fu_8559_p1 == 10'd243) & ~(trunc_ln321_fu_8559_p1 == 10'd242) & ~(trunc_ln321_fu_8559_p1 == 10'd241) & ~(trunc_ln321_fu_8559_p1 == 10'd240) & ~(trunc_ln321_fu_8559_p1 == 10'd239) & ~(trunc_ln321_fu_8559_p1 == 10'd238) & ~(trunc_ln321_fu_8559_p1 == 10'd237) & ~(trunc_ln321_fu_8559_p1 == 10'd236) & ~(trunc_ln321_fu_8559_p1 == 10'd235) & ~(trunc_ln321_fu_8559_p1 == 10'd234) & ~(trunc_ln321_fu_8559_p1 == 10'd233) & ~(trunc_ln321_fu_8559_p1 == 10'd232) & ~(trunc_ln321_fu_8559_p1 == 10'd231) & ~(trunc_ln321_fu_8559_p1 == 10'd230) & ~(trunc_ln321_fu_8559_p1 == 10'd229) & ~(trunc_ln321_fu_8559_p1 == 10'd228) & ~(trunc_ln321_fu_8559_p1 == 10'd227) & ~(trunc_ln321_fu_8559_p1 == 10'd226) & ~(trunc_ln321_fu_8559_p1 == 10'd225) & ~(trunc_ln321_fu_8559_p1 == 10'd224) & ~(trunc_ln321_fu_8559_p1 == 10'd223) & ~(trunc_ln321_fu_8559_p1 == 10'd222) & ~(trunc_ln321_fu_8559_p1 == 10'd221) & ~(trunc_ln321_fu_8559_p1 == 10'd220) & ~(trunc_ln321_fu_8559_p1 == 10'd219) & ~(trunc_ln321_fu_8559_p1 == 10'd218) & ~(trunc_ln321_fu_8559_p1 == 10'd217) & ~(trunc_ln321_fu_8559_p1 == 10'd216) & ~(trunc_ln321_fu_8559_p1 == 10'd215) & ~(trunc_ln321_fu_8559_p1 == 10'd214) & ~(trunc_ln321_fu_8559_p1 == 10'd213) & ~(trunc_ln321_fu_8559_p1 == 10'd212) & ~(trunc_ln321_fu_8559_p1 == 10'd211) & ~(trunc_ln321_fu_8559_p1 == 10'd210) & ~(trunc_ln321_fu_8559_p1 == 10'd209) & ~(trunc_ln321_fu_8559_p1 == 10'd208) & ~(trunc_ln321_fu_8559_p1 == 10'd207) & ~(trunc_ln321_fu_8559_p1 == 10'd206) & ~(trunc_ln321_fu_8559_p1 == 10'd205) & ~(trunc_ln321_fu_8559_p1 == 10'd204) & ~(trunc_ln321_fu_8559_p1 == 10'd203) & ~(trunc_ln321_fu_8559_p1 == 10'd202) & ~(trunc_ln321_fu_8559_p1 == 10'd201) & ~(trunc_ln321_fu_8559_p1 == 10'd200) & ~(trunc_ln321_fu_8559_p1 == 10'd199) & ~(trunc_ln321_fu_8559_p1 == 10'd198) & ~(trunc_ln321_fu_8559_p1 == 10'd197) & ~(trunc_ln321_fu_8559_p1 == 10'd196) & ~(trunc_ln321_fu_8559_p1 == 10'd195) & ~(trunc_ln321_fu_8559_p1 == 10'd194) & ~(trunc_ln321_fu_8559_p1 == 10'd193) & ~(trunc_ln321_fu_8559_p1 == 10'd192) & ~(trunc_ln321_fu_8559_p1 == 10'd191) & ~(trunc_ln321_fu_8559_p1 == 10'd190) & ~(trunc_ln321_fu_8559_p1 == 10'd189) & ~(trunc_ln321_fu_8559_p1 == 10'd188) & ~(trunc_ln321_fu_8559_p1 == 10'd187) & ~(trunc_ln321_fu_8559_p1 == 10'd186) & ~(trunc_ln321_fu_8559_p1 == 10'd185) & ~(trunc_ln321_fu_8559_p1 == 10'd184) & ~(trunc_ln321_fu_8559_p1 == 10'd183) & ~(trunc_ln321_fu_8559_p1 == 10'd182) & ~(trunc_ln321_fu_8559_p1 == 10'd181) & ~(trunc_ln321_fu_8559_p1 == 10'd180) & ~(trunc_ln321_fu_8559_p1 == 10'd179) & ~(trunc_ln321_fu_8559_p1 == 10'd178) & ~(trunc_ln321_fu_8559_p1 == 10'd177) & ~(trunc_ln321_fu_8559_p1 == 10'd176) & ~(trunc_ln321_fu_8559_p1 == 10'd175) & ~(trunc_ln321_fu_8559_p1 == 10'd174) & ~(trunc_ln321_fu_8559_p1 == 10'd173) & ~(trunc_ln321_fu_8559_p1 == 10'd172) & ~(trunc_ln321_fu_8559_p1 == 10'd171) & ~(trunc_ln321_fu_8559_p1 == 10'd170) & ~(trunc_ln321_fu_8559_p1 == 10'd169) & ~(trunc_ln321_fu_8559_p1 == 10'd168) & ~(trunc_ln321_fu_8559_p1 == 10'd167) & ~(trunc_ln321_fu_8559_p1 == 10'd166) & ~(trunc_ln321_fu_8559_p1 == 10'd165) & ~(trunc_ln321_fu_8559_p1 == 10'd164) & ~(trunc_ln321_fu_8559_p1 == 10'd163) & ~(trunc_ln321_fu_8559_p1 == 10'd162) & ~(trunc_ln321_fu_8559_p1 == 10'd161) & ~(trunc_ln321_fu_8559_p1 == 10'd160) & ~(trunc_ln321_fu_8559_p1 == 10'd159) & ~(trunc_ln321_fu_8559_p1 == 10'd158) & ~(trunc_ln321_fu_8559_p1 == 10'd157) & ~(trunc_ln321_fu_8559_p1 == 10'd156) & ~(trunc_ln321_fu_8559_p1 == 10'd155) & ~(trunc_ln321_fu_8559_p1 == 10'd154) & ~(trunc_ln321_fu_8559_p1 == 10'd153) & ~(trunc_ln321_fu_8559_p1 == 10'd152) & ~(trunc_ln321_fu_8559_p1 == 10'd151) & ~(trunc_ln321_fu_8559_p1 == 10'd150) & ~(trunc_ln321_fu_8559_p1 == 10'd149) & ~(trunc_ln321_fu_8559_p1 == 10'd148) & ~(trunc_ln321_fu_8559_p1 == 10'd147) & ~(trunc_ln321_fu_8559_p1 == 10'd146) & ~(trunc_ln321_fu_8559_p1 == 10'd145) & ~(trunc_ln321_fu_8559_p1 == 10'd144) & ~(trunc_ln321_fu_8559_p1 == 10'd143) & ~(trunc_ln321_fu_8559_p1 == 10'd142) & ~(trunc_ln321_fu_8559_p1 == 10'd141) & ~(trunc_ln321_fu_8559_p1 == 10'd140) & ~(trunc_ln321_fu_8559_p1 == 10'd139) & ~(trunc_ln321_fu_8559_p1 == 10'd138) & ~(trunc_ln321_fu_8559_p1 == 10'd137) & ~(trunc_ln321_fu_8559_p1 == 10'd136) & ~(trunc_ln321_fu_8559_p1 == 10'd135) & ~(trunc_ln321_fu_8559_p1 == 10'd134) & ~(trunc_ln321_fu_8559_p1 == 10'd133) & ~(trunc_ln321_fu_8559_p1 == 10'd132) & ~(trunc_ln321_fu_8559_p1 == 10'd131) & ~(trunc_ln321_fu_8559_p1 == 10'd130) & ~(trunc_ln321_fu_8559_p1 == 10'd129) & ~(trunc_ln321_fu_8559_p1 == 10'd128) & ~(trunc_ln321_fu_8559_p1 == 10'd127) & ~(trunc_ln321_fu_8559_p1 == 10'd126) & ~(trunc_ln321_fu_8559_p1 == 10'd125) & ~(trunc_ln321_fu_8559_p1 == 10'd124) & ~(trunc_ln321_fu_8559_p1 == 10'd123) & ~(trunc_ln321_fu_8559_p1 == 10'd122) & ~(trunc_ln321_fu_8559_p1 == 10'd121) & ~(trunc_ln321_fu_8559_p1 == 10'd120) & ~(trunc_ln321_fu_8559_p1 == 10'd119) & ~(trunc_ln321_fu_8559_p1 == 10'd118) & ~(trunc_ln321_fu_8559_p1 == 10'd117) & ~(trunc_ln321_fu_8559_p1 == 10'd116) & ~(trunc_ln321_fu_8559_p1 == 10'd115) & ~(trunc_ln321_fu_8559_p1 == 10'd114) & ~(trunc_ln321_fu_8559_p1 == 10'd113) & ~(trunc_ln321_fu_8559_p1 == 10'd112) & ~(trunc_ln321_fu_8559_p1 == 10'd111) & ~(trunc_ln321_fu_8559_p1 == 10'd110) & ~(trunc_ln321_fu_8559_p1 == 10'd109) & ~(trunc_ln321_fu_8559_p1 == 10'd108) & ~(trunc_ln321_fu_8559_p1 == 10'd107) & ~(trunc_ln321_fu_8559_p1 == 10'd106) & ~(trunc_ln321_fu_8559_p1 == 10'd105) & ~(trunc_ln321_fu_8559_p1 == 10'd104) & ~(trunc_ln321_fu_8559_p1 == 10'd103) & ~(trunc_ln321_fu_8559_p1 == 10'd102) & ~(trunc_ln321_fu_8559_p1 == 10'd101) & ~(trunc_ln321_fu_8559_p1 == 10'd100) & ~(trunc_ln321_fu_8559_p1 == 10'd99) & ~(trunc_ln321_fu_8559_p1 == 10'd98) & ~(trunc_ln321_fu_8559_p1 == 10'd97) & ~(trunc_ln321_fu_8559_p1 == 10'd96) & ~(trunc_ln321_fu_8559_p1 == 10'd95) & ~(trunc_ln321_fu_8559_p1 == 10'd94) & ~(trunc_ln321_fu_8559_p1 == 10'd93) & ~(trunc_ln321_fu_8559_p1 == 10'd92) & ~(trunc_ln321_fu_8559_p1 == 10'd91) & ~(trunc_ln321_fu_8559_p1 == 10'd90) & ~(trunc_ln321_fu_8559_p1 == 10'd89) & ~(trunc_ln321_fu_8559_p1 == 10'd88) & ~(trunc_ln321_fu_8559_p1 == 10'd87) & ~(trunc_ln321_fu_8559_p1 == 10'd86) & ~(trunc_ln321_fu_8559_p1 == 10'd85) & ~(trunc_ln321_fu_8559_p1 == 10'd84) & ~(trunc_ln321_fu_8559_p1 == 10'd83) & ~(trunc_ln321_fu_8559_p1 == 10'd82) & ~(trunc_ln321_fu_8559_p1 == 10'd81) & ~(trunc_ln321_fu_8559_p1 == 10'd80) & ~(trunc_ln321_fu_8559_p1 == 10'd79) & ~(trunc_ln321_fu_8559_p1 == 10'd78) & ~(trunc_ln321_fu_8559_p1 == 10'd77) & ~(trunc_ln321_fu_8559_p1 == 10'd76) & ~(trunc_ln321_fu_8559_p1 == 10'd75) & ~(trunc_ln321_fu_8559_p1 == 10'd74) & ~(trunc_ln321_fu_8559_p1 == 10'd73) & ~(trunc_ln321_fu_8559_p1 == 10'd72) & ~(trunc_ln321_fu_8559_p1 == 10'd71) & ~(trunc_ln321_fu_8559_p1 == 10'd70) & ~(trunc_ln321_fu_8559_p1 == 10'd69) & ~(trunc_ln321_fu_8559_p1 == 10'd68) & ~(trunc_ln321_fu_8559_p1 == 10'd67) & ~(trunc_ln321_fu_8559_p1 == 10'd66) & ~(trunc_ln321_fu_8559_p1 == 10'd65) & ~(trunc_ln321_fu_8559_p1 == 10'd64) & ~(trunc_ln321_fu_8559_p1 == 10'd63) & ~(trunc_ln321_fu_8559_p1 == 10'd62) & ~(trunc_ln321_fu_8559_p1 == 10'd61) & ~(trunc_ln321_fu_8559_p1 == 10'd60) & ~(trunc_ln321_fu_8559_p1 == 10'd59) & ~(trunc_ln321_fu_8559_p1 == 10'd58) & ~(trunc_ln321_fu_8559_p1 == 10'd57) & ~(trunc_ln321_fu_8559_p1 == 10'd56) & ~(trunc_ln321_fu_8559_p1 == 10'd55) & ~(trunc_ln321_fu_8559_p1 == 10'd54) & ~(trunc_ln321_fu_8559_p1 == 10'd53) & ~(trunc_ln321_fu_8559_p1 == 10'd52) & ~(trunc_ln321_fu_8559_p1 == 10'd51) & ~(trunc_ln321_fu_8559_p1 == 10'd50) & ~(trunc_ln321_fu_8559_p1 == 10'd49) & ~(trunc_ln321_fu_8559_p1 == 10'd48) & ~(trunc_ln321_fu_8559_p1 == 10'd47) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_576_fu_3710 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd56) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_57_fu_1634 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd57) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_58_fu_1638 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd58) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_59_fu_1642 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd4) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_5_fu_1426 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd59) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_60_fu_1646 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd60) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_61_fu_1650 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd61) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_62_fu_1654 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd62) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_63_fu_1658 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd63) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_64_fu_1662 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd64) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_65_fu_1666 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd65) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_66_fu_1670 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd66) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_67_fu_1674 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd67) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_68_fu_1678 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd68) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_69_fu_1682 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd5) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_6_fu_1430 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd69) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_70_fu_1686 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd70) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_71_fu_1690 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd71) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_72_fu_1694 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd72) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_73_fu_1698 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd73) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_74_fu_1702 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd74) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_75_fu_1706 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd75) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_76_fu_1710 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd76) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_77_fu_1714 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd77) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_78_fu_1718 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd78) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_79_fu_1722 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd6) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_7_fu_1434 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd79) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_80_fu_1726 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd80) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_81_fu_1730 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd81) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_82_fu_1734 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd82) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_83_fu_1738 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd83) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_84_fu_1742 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd84) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_85_fu_1746 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd85) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_86_fu_1750 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd86) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_87_fu_1754 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd87) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_88_fu_1758 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd88) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_89_fu_1762 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd7) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_8_fu_1438 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd89) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_90_fu_1766 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd90) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_91_fu_1770 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd91) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_92_fu_1774 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd92) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_93_fu_1778 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd93) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_94_fu_1782 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd94) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_95_fu_1786 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd95) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_96_fu_1790 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd96) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_97_fu_1794 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd97) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_98_fu_1798 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd98) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_99_fu_1802 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd8) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_9_fu_1442 <= in_V_V_TDATA;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln321_fu_8559_p1 == 10'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_V_fu_1410 <= in_V_V_TDATA;
    end
end

always @ (*) begin
    if ((icmp_ln248_fu_5645_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state6) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_17768 == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_sig_allocacmp_nf_assign_load_1 = select_ln301_fu_11988_p3;
    end else begin
        ap_sig_allocacmp_nf_assign_load_1 = nf_assign_fu_3714;
    end
end

always @ (*) begin
    if (((icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_predicate_op1185_read_state2 == 1'b1))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln289_reg_17768_pp0_iter2_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln289_reg_17768_pp0_iter2_reg == 1'd1) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_10_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_10_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_11_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_11_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_12_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_12_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_13_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_13_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_14_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_14_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_15_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_15_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_16_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_16_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_17_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_17_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_18_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_18_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_19_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_19_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_1_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_1_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_20_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_20_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_21_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_21_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_22_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_22_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_23_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_23_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_24_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_24_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_25_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_25_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_26_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_26_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_27_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_27_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_28_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_28_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_29_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_29_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_2_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_2_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_30_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_30_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_31_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_31_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_32_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_32_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_33_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_33_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_34_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_34_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_35_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_35_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_36_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_36_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_37_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_37_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_38_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_38_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_39_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_39_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_3_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_3_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_40_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_40_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_41_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_41_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_42_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_42_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_43_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_43_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_44_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_44_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_45_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_45_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_46_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_46_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_47_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_47_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_48_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_48_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_49_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_49_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_4_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_4_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_50_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_50_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_51_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_51_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_52_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_52_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_53_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_53_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_54_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_54_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_55_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_55_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_5_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_5_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_6_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_6_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_7_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_7_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_8_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_8_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_9_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_9_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        threshs_m_thresholds_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln248_fu_5645_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TDATA_blk_n = weight_V_V_TVALID;
    end else begin
        weight_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln248_fu_5645_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_V_V_TREADY = 1'b1;
    end else begin
        weight_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln248_fu_5645_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((ap_enable_reg_pp0_iter2 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter2 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (icmp_ln248_fu_5645_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accu_0_0_V_fu_12053_p2 = ($signed(add_ln700_fu_12044_p2) + $signed(sext_ln700_2_fu_12050_p1));

assign accu_0_1_V_fu_12071_p2 = ($signed(add_ln700_4_fu_12062_p2) + $signed(sext_ln700_5_fu_12068_p1));

assign accu_0_2_V_fu_12089_p2 = ($signed(add_ln700_8_fu_12080_p2) + $signed(sext_ln700_8_fu_12086_p1));

assign accu_0_3_V_fu_12107_p2 = ($signed(add_ln700_12_fu_12098_p2) + $signed(sext_ln700_11_fu_12104_p1));

assign add_ln700_10_fu_11847_p2 = ($signed(sext_ln170_5_fu_11824_p1) + $signed(add_ln700_9_fu_11841_p2));

assign add_ln700_12_fu_12098_p2 = ($signed(sext_ln700_9_fu_12095_p1) + $signed(select_ln271_fu_12013_p3));

assign add_ln700_13_fu_11901_p2 = ($signed(sext_ln700_10_fu_11897_p1) + $signed(sext_ln170_6_fu_11862_p1));

assign add_ln700_14_fu_11907_p2 = ($signed(sext_ln170_7_fu_11884_p1) + $signed(add_ln700_13_fu_11901_p2));

assign add_ln700_16_fu_12751_p2 = (zext_ln142_2_fu_12639_p1 + zext_ln142_3_fu_12648_p1);

assign add_ln700_17_fu_12757_p2 = (add_ln700_16_fu_12751_p2 + zext_ln142_1_fu_12630_p1);

assign add_ln700_18_fu_12767_p2 = (zext_ln142_4_fu_12657_p1 + zext_ln142_5_fu_12666_p1);

assign add_ln700_19_fu_12777_p2 = (zext_ln142_6_fu_12675_p1 + zext_ln142_7_fu_12684_p1);

assign add_ln700_1_fu_11721_p2 = ($signed(sext_ln700_1_fu_11717_p1) + $signed(sext_ln170_fu_11640_p1));

assign add_ln700_20_fu_12787_p2 = (zext_ln700_3_fu_12783_p1 + zext_ln700_2_fu_12773_p1);

assign add_ln700_21_fu_12793_p2 = (add_ln700_20_fu_12787_p2 + zext_ln700_1_fu_12763_p1);

assign add_ln700_22_fu_12803_p2 = (zext_ln142_9_fu_12702_p1 + zext_ln142_10_fu_12711_p1);

assign add_ln700_23_fu_12809_p2 = (add_ln700_22_fu_12803_p2 + zext_ln142_8_fu_12693_p1);

assign add_ln700_24_fu_12819_p2 = (zext_ln142_11_fu_12720_p1 + zext_ln142_12_fu_12729_p1);

assign add_ln700_25_fu_12829_p2 = (zext_ln142_13_fu_12738_p1 + zext_ln700_fu_12747_p1);

assign add_ln700_26_fu_12839_p2 = (zext_ln700_7_fu_12835_p1 + zext_ln700_6_fu_12825_p1);

assign add_ln700_27_fu_12845_p2 = (add_ln700_26_fu_12839_p2 + zext_ln700_5_fu_12815_p1);

assign add_ln700_28_fu_12855_p2 = (zext_ln700_8_fu_12851_p1 + zext_ln700_4_fu_12799_p1);

assign add_ln700_29_fu_12987_p2 = (zext_ln142_15_fu_12875_p1 + zext_ln142_16_fu_12884_p1);

assign add_ln700_2_fu_11727_p2 = ($signed(sext_ln170_1_fu_11690_p1) + $signed(add_ln700_1_fu_11721_p2));

assign add_ln700_30_fu_12993_p2 = (add_ln700_29_fu_12987_p2 + zext_ln142_14_fu_12866_p1);

assign add_ln700_31_fu_13003_p2 = (zext_ln142_17_fu_12893_p1 + zext_ln142_18_fu_12902_p1);

assign add_ln700_32_fu_13013_p2 = (zext_ln142_19_fu_12911_p1 + zext_ln142_20_fu_12920_p1);

assign add_ln700_33_fu_13023_p2 = (zext_ln700_12_fu_13019_p1 + zext_ln700_11_fu_13009_p1);

assign add_ln700_34_fu_13029_p2 = (add_ln700_33_fu_13023_p2 + zext_ln700_10_fu_12999_p1);

assign add_ln700_35_fu_13039_p2 = (zext_ln142_22_fu_12938_p1 + zext_ln142_23_fu_12947_p1);

assign add_ln700_36_fu_13045_p2 = (add_ln700_35_fu_13039_p2 + zext_ln142_21_fu_12929_p1);

assign add_ln700_37_fu_13055_p2 = (zext_ln142_24_fu_12956_p1 + zext_ln142_25_fu_12965_p1);

assign add_ln700_38_fu_13065_p2 = (zext_ln142_26_fu_12974_p1 + zext_ln700_9_fu_12983_p1);

assign add_ln700_39_fu_13075_p2 = (zext_ln700_16_fu_13071_p1 + zext_ln700_15_fu_13061_p1);

assign add_ln700_40_fu_13081_p2 = (add_ln700_39_fu_13075_p2 + zext_ln700_14_fu_13051_p1);

assign add_ln700_41_fu_13091_p2 = (zext_ln700_17_fu_13087_p1 + zext_ln700_13_fu_13035_p1);

assign add_ln700_42_fu_13223_p2 = (zext_ln142_28_fu_13111_p1 + zext_ln142_29_fu_13120_p1);

assign add_ln700_43_fu_13229_p2 = (add_ln700_42_fu_13223_p2 + zext_ln142_27_fu_13102_p1);

assign add_ln700_44_fu_13239_p2 = (zext_ln142_30_fu_13129_p1 + zext_ln142_31_fu_13138_p1);

assign add_ln700_45_fu_13249_p2 = (zext_ln142_32_fu_13147_p1 + zext_ln142_33_fu_13156_p1);

assign add_ln700_46_fu_13259_p2 = (zext_ln700_21_fu_13255_p1 + zext_ln700_20_fu_13245_p1);

assign add_ln700_47_fu_13265_p2 = (add_ln700_46_fu_13259_p2 + zext_ln700_19_fu_13235_p1);

assign add_ln700_48_fu_13275_p2 = (zext_ln142_35_fu_13174_p1 + zext_ln142_36_fu_13183_p1);

assign add_ln700_49_fu_13281_p2 = (add_ln700_48_fu_13275_p2 + zext_ln142_34_fu_13165_p1);

assign add_ln700_4_fu_12062_p2 = ($signed(sext_ln700_3_fu_12059_p1) + $signed(select_ln271_2_fu_12027_p3));

assign add_ln700_50_fu_13291_p2 = (zext_ln142_37_fu_13192_p1 + zext_ln142_38_fu_13201_p1);

assign add_ln700_51_fu_13301_p2 = (zext_ln142_39_fu_13210_p1 + zext_ln700_18_fu_13219_p1);

assign add_ln700_52_fu_13311_p2 = (zext_ln700_25_fu_13307_p1 + zext_ln700_24_fu_13297_p1);

assign add_ln700_53_fu_13317_p2 = (add_ln700_52_fu_13311_p2 + zext_ln700_23_fu_13287_p1);

assign add_ln700_54_fu_13327_p2 = (zext_ln700_26_fu_13323_p1 + zext_ln700_22_fu_13271_p1);

assign add_ln700_55_fu_13459_p2 = (zext_ln142_41_fu_13347_p1 + zext_ln142_42_fu_13356_p1);

assign add_ln700_56_fu_13465_p2 = (add_ln700_55_fu_13459_p2 + zext_ln142_40_fu_13338_p1);

assign add_ln700_57_fu_13475_p2 = (zext_ln142_43_fu_13365_p1 + zext_ln142_44_fu_13374_p1);

assign add_ln700_58_fu_13485_p2 = (zext_ln142_45_fu_13383_p1 + zext_ln142_46_fu_13392_p1);

assign add_ln700_59_fu_13495_p2 = (zext_ln700_30_fu_13491_p1 + zext_ln700_29_fu_13481_p1);

assign add_ln700_5_fu_11781_p2 = ($signed(sext_ln700_4_fu_11777_p1) + $signed(sext_ln170_2_fu_11742_p1));

assign add_ln700_60_fu_13501_p2 = (add_ln700_59_fu_13495_p2 + zext_ln700_28_fu_13471_p1);

assign add_ln700_61_fu_13511_p2 = (zext_ln142_48_fu_13410_p1 + zext_ln142_49_fu_13419_p1);

assign add_ln700_62_fu_13517_p2 = (add_ln700_61_fu_13511_p2 + zext_ln142_47_fu_13401_p1);

assign add_ln700_63_fu_13527_p2 = (zext_ln142_50_fu_13428_p1 + zext_ln142_51_fu_13437_p1);

assign add_ln700_64_fu_13537_p2 = (zext_ln142_52_fu_13446_p1 + zext_ln700_27_fu_13455_p1);

assign add_ln700_65_fu_13547_p2 = (zext_ln700_34_fu_13543_p1 + zext_ln700_33_fu_13533_p1);

assign add_ln700_66_fu_13553_p2 = (add_ln700_65_fu_13547_p2 + zext_ln700_32_fu_13523_p1);

assign add_ln700_67_fu_13563_p2 = (zext_ln700_35_fu_13559_p1 + zext_ln700_31_fu_13507_p1);

assign add_ln700_6_fu_11787_p2 = ($signed(sext_ln170_3_fu_11764_p1) + $signed(add_ln700_5_fu_11781_p2));

assign add_ln700_8_fu_12080_p2 = ($signed(sext_ln700_6_fu_12077_p1) + $signed(select_ln271_1_fu_12020_p3));

assign add_ln700_9_fu_11841_p2 = ($signed(sext_ln700_7_fu_11837_p1) + $signed(sext_ln170_4_fu_11802_p1));

assign add_ln700_fu_12044_p2 = ($signed(sext_ln700_fu_12041_p1) + $signed(select_ln271_3_fu_12034_p3));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state6 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op1185_read_state2 == 1'b1)) | ((icmp_ln248_fu_5645_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_block_state5_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op1185_read_state2 == 1'b1)) | ((icmp_ln248_fu_5645_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_block_state5_io)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (((in_V_V_TVALID == 1'b0) & (ap_predicate_op1185_read_state2 == 1'b1)) | ((icmp_ln248_fu_5645_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)))));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = (((in_V_V_TVALID == 1'b0) & (ap_predicate_op1185_read_state2 == 1'b1)) | ((icmp_ln248_fu_5645_p2 == 1'd0) & (weight_V_V_TVALID == 1'b0)));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state5_io = ((icmp_ln289_reg_17768_pp0_iter2_reg == 1'd1) & (out_V_V_TREADY == 1'b0));
end

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_reg_pp0_iter0_act_m_val_V_reg_4476 = 'bx;

always @ (*) begin
    ap_predicate_op1185_read_state2 = ((icmp_ln252_fu_5660_p2 == 1'd1) & (icmp_ln248_fu_5645_p2 == 1'd0));
end

assign arg_V_read_assign_1_fu_11644_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_4476[7:4]}};

assign arg_V_read_assign_2_fu_11667_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_4476[11:8]}};

assign arg_V_read_assign_3_fu_11694_p4 = {{ap_phi_reg_pp0_iter1_act_m_val_V_reg_4476[15:12]}};

assign i_fu_5651_p2 = (i_0_reg_4465 + 16'd1);

assign icmp_ln248_fu_5645_p2 = ((i_0_reg_4465 == 16'd36864) ? 1'b1 : 1'b0);

assign icmp_ln252_fu_5660_p2 = ((ap_sig_allocacmp_nf_assign_load_1 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln271_fu_11446_p2 = ((sf_1_fu_1406 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln289_fu_11612_p2 = ((sf_fu_11606_p2 == 32'd576) ? 1'b1 : 1'b0);

assign icmp_ln301_fu_11982_p2 = ((nf_fu_11976_p2 == 32'd64) ? 1'b1 : 1'b0);

assign icmp_ln899_10_fu_12237_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_10_fu_12233_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_11_fu_12247_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_11_fu_12243_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_12_fu_12257_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_12_fu_12253_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_13_fu_12267_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_13_fu_12263_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_14_fu_12273_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_41_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_15_fu_12279_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_40_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_16_fu_12285_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_35_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_17_fu_12291_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_34_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_18_fu_12297_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_33_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_19_fu_12303_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_32_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_1_fu_12147_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_1_fu_12143_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_20_fu_12309_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_31_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_21_fu_12315_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_30_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_22_fu_12321_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_29_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_23_fu_12327_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_28_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_24_fu_12333_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_39_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_25_fu_12339_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_38_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_26_fu_12345_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_37_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_27_fu_12351_p2 = (($signed(accu_0_1_V_fu_12071_p2) < $signed(threshs_m_thresholds_36_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_28_fu_12361_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_14_fu_12357_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_29_fu_12371_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_15_fu_12367_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_2_fu_12157_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_2_fu_12153_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_30_fu_12381_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_16_fu_12377_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_31_fu_12391_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_17_fu_12387_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_32_fu_12401_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_18_fu_12397_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_33_fu_12411_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_19_fu_12407_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_34_fu_12421_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_20_fu_12417_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_35_fu_12431_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_21_fu_12427_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_36_fu_12441_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_22_fu_12437_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_37_fu_12451_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_23_fu_12447_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_38_fu_12461_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_24_fu_12457_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_39_fu_12471_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_25_fu_12467_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_3_fu_12167_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_3_fu_12163_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_40_fu_12481_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_26_fu_12477_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_41_fu_12491_p2 = (($signed(accu_0_2_V_fu_12089_p2) < $signed(sext_ln142_27_fu_12487_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_42_fu_12497_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(threshs_m_thresholds_13_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_43_fu_12507_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_28_fu_12503_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_44_fu_12517_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_29_fu_12513_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_45_fu_12527_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_30_fu_12523_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_46_fu_12537_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_31_fu_12533_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_47_fu_12547_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_32_fu_12543_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_48_fu_12557_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_33_fu_12553_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_49_fu_12567_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_34_fu_12563_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_4_fu_12177_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_4_fu_12173_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_50_fu_12577_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_35_fu_12573_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_51_fu_12587_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_36_fu_12583_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_52_fu_12597_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_37_fu_12593_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_53_fu_12607_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(sext_ln142_38_fu_12603_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_54_fu_12613_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(threshs_m_thresholds_9_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_55_fu_12619_p2 = (($signed(accu_0_3_V_fu_12107_p2) < $signed(threshs_m_thresholds_8_q0)) ? 1'b1 : 1'b0);

assign icmp_ln899_5_fu_12187_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_5_fu_12183_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_6_fu_12197_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_6_fu_12193_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_7_fu_12207_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_7_fu_12203_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_8_fu_12217_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_8_fu_12213_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_9_fu_12227_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_9_fu_12223_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_fu_12137_p2 = (($signed(accu_0_0_V_fu_12053_p2) < $signed(sext_ln142_fu_12133_p1)) ? 1'b1 : 1'b0);

assign inElem_V_1_fu_7401_p577 = sf_1_fu_1406[9:0];

assign mul_ln1352_10_fu_11818_p0 = sext_ln215_5_fu_11680_p1;

assign mul_ln1352_11_fu_11831_p0 = sext_ln215_7_fu_11707_p1;

assign mul_ln1352_12_fu_11856_p0 = sext_ln215_1_fu_11630_p1;

assign mul_ln1352_13_fu_11869_p0 = sext_ln215_3_fu_11657_p1;

assign mul_ln1352_14_fu_11878_p0 = sext_ln215_5_fu_11680_p1;

assign mul_ln1352_15_fu_11891_p0 = sext_ln215_7_fu_11707_p1;

assign mul_ln1352_1_fu_11661_p0 = sext_ln215_3_fu_11657_p1;

assign mul_ln1352_2_fu_11684_p0 = sext_ln215_5_fu_11680_p1;

assign mul_ln1352_3_fu_11711_p0 = sext_ln215_7_fu_11707_p1;

assign mul_ln1352_4_fu_11736_p0 = sext_ln215_1_fu_11630_p1;

assign mul_ln1352_5_fu_11749_p0 = sext_ln215_3_fu_11657_p1;

assign mul_ln1352_6_fu_11758_p0 = sext_ln215_5_fu_11680_p1;

assign mul_ln1352_7_fu_11771_p0 = sext_ln215_7_fu_11707_p1;

assign mul_ln1352_8_fu_11796_p0 = sext_ln215_1_fu_11630_p1;

assign mul_ln1352_9_fu_11809_p0 = sext_ln215_3_fu_11657_p1;

assign mul_ln1352_fu_11634_p0 = sext_ln215_1_fu_11630_p1;

assign nf_fu_11976_p2 = (nf_assign_fu_3714 + 32'd1);

assign out_V_V_TDATA = {{{{add_ln700_67_fu_13563_p2}, {add_ln700_54_fu_13327_p2}}, {add_ln700_41_fu_13091_p2}}, {add_ln700_28_fu_12855_p2}};

assign select_ln271_1_fu_12020_p3 = ((icmp_ln271_reg_17680_pp0_iter1_reg[0:0] === 1'b1) ? 18'd0 : accu_V_0_2_0_fu_1398);

assign select_ln271_2_fu_12027_p3 = ((icmp_ln271_reg_17680_pp0_iter1_reg[0:0] === 1'b1) ? 18'd0 : accu_V_0_1_0_fu_1394);

assign select_ln271_3_fu_12034_p3 = ((icmp_ln271_reg_17680_pp0_iter1_reg[0:0] === 1'b1) ? 18'd0 : accu_V_0_0_0_fu_1390);

assign select_ln271_fu_12013_p3 = ((icmp_ln271_reg_17680_pp0_iter1_reg[0:0] === 1'b1) ? 18'd0 : accu_V_0_3_0_fu_1402);

assign select_ln301_fu_11988_p3 = ((icmp_ln301_fu_11982_p2[0:0] === 1'b1) ? 32'd0 : nf_fu_11976_p2);

assign sext_ln142_10_fu_12233_p1 = $signed(threshs_m_thresholds_53_q0);

assign sext_ln142_11_fu_12243_p1 = $signed(threshs_m_thresholds_52_q0);

assign sext_ln142_12_fu_12253_p1 = $signed(threshs_m_thresholds_51_q0);

assign sext_ln142_13_fu_12263_p1 = $signed(threshs_m_thresholds_50_q0);

assign sext_ln142_14_fu_12357_p1 = $signed(threshs_m_thresholds_27_q0);

assign sext_ln142_15_fu_12367_p1 = $signed(threshs_m_thresholds_26_q0);

assign sext_ln142_16_fu_12377_p1 = $signed(threshs_m_thresholds_21_q0);

assign sext_ln142_17_fu_12387_p1 = $signed(threshs_m_thresholds_20_q0);

assign sext_ln142_18_fu_12397_p1 = $signed(threshs_m_thresholds_19_q0);

assign sext_ln142_19_fu_12407_p1 = $signed(threshs_m_thresholds_18_q0);

assign sext_ln142_1_fu_12143_p1 = $signed(threshs_m_thresholds_54_q0);

assign sext_ln142_20_fu_12417_p1 = $signed(threshs_m_thresholds_17_q0);

assign sext_ln142_21_fu_12427_p1 = $signed(threshs_m_thresholds_16_q0);

assign sext_ln142_22_fu_12437_p1 = $signed(threshs_m_thresholds_15_q0);

assign sext_ln142_23_fu_12447_p1 = $signed(threshs_m_thresholds_14_q0);

assign sext_ln142_24_fu_12457_p1 = $signed(threshs_m_thresholds_25_q0);

assign sext_ln142_25_fu_12467_p1 = $signed(threshs_m_thresholds_24_q0);

assign sext_ln142_26_fu_12477_p1 = $signed(threshs_m_thresholds_23_q0);

assign sext_ln142_27_fu_12487_p1 = $signed(threshs_m_thresholds_22_q0);

assign sext_ln142_28_fu_12503_p1 = $signed(threshs_m_thresholds_12_q0);

assign sext_ln142_29_fu_12513_p1 = $signed(threshs_m_thresholds_7_q0);

assign sext_ln142_2_fu_12153_p1 = $signed(threshs_m_thresholds_49_q0);

assign sext_ln142_30_fu_12523_p1 = $signed(threshs_m_thresholds_6_q0);

assign sext_ln142_31_fu_12533_p1 = $signed(threshs_m_thresholds_5_q0);

assign sext_ln142_32_fu_12543_p1 = $signed(threshs_m_thresholds_4_q0);

assign sext_ln142_33_fu_12553_p1 = $signed(threshs_m_thresholds_3_q0);

assign sext_ln142_34_fu_12563_p1 = $signed(threshs_m_thresholds_2_q0);

assign sext_ln142_35_fu_12573_p1 = $signed(threshs_m_thresholds_1_q0);

assign sext_ln142_36_fu_12583_p1 = $signed(threshs_m_thresholds_q0);

assign sext_ln142_37_fu_12593_p1 = $signed(threshs_m_thresholds_11_q0);

assign sext_ln142_38_fu_12603_p1 = $signed(threshs_m_thresholds_10_q0);

assign sext_ln142_3_fu_12163_p1 = $signed(threshs_m_thresholds_48_q0);

assign sext_ln142_4_fu_12173_p1 = $signed(threshs_m_thresholds_47_q0);

assign sext_ln142_5_fu_12183_p1 = $signed(threshs_m_thresholds_46_q0);

assign sext_ln142_6_fu_12193_p1 = $signed(threshs_m_thresholds_45_q0);

assign sext_ln142_7_fu_12203_p1 = $signed(threshs_m_thresholds_44_q0);

assign sext_ln142_8_fu_12213_p1 = $signed(threshs_m_thresholds_43_q0);

assign sext_ln142_9_fu_12223_p1 = $signed(threshs_m_thresholds_42_q0);

assign sext_ln142_fu_12133_p1 = $signed(threshs_m_thresholds_55_q0);

assign sext_ln170_1_fu_11690_p1 = mul_ln1352_2_fu_11684_p2;

assign sext_ln170_2_fu_11742_p1 = mul_ln1352_4_fu_11736_p2;

assign sext_ln170_3_fu_11764_p1 = mul_ln1352_6_fu_11758_p2;

assign sext_ln170_4_fu_11802_p1 = mul_ln1352_8_fu_11796_p2;

assign sext_ln170_5_fu_11824_p1 = mul_ln1352_10_fu_11818_p2;

assign sext_ln170_6_fu_11862_p1 = mul_ln1352_12_fu_11856_p2;

assign sext_ln170_7_fu_11884_p1 = mul_ln1352_14_fu_11878_p2;

assign sext_ln170_fu_11640_p1 = mul_ln1352_fu_11634_p2;

assign sext_ln215_1_fu_11630_p1 = $signed(trunc_ln647_1_fu_11623_p1);

assign sext_ln215_3_fu_11657_p1 = $signed(arg_V_read_assign_1_fu_11644_p4);

assign sext_ln215_5_fu_11680_p1 = $signed(arg_V_read_assign_2_fu_11667_p4);

assign sext_ln215_7_fu_11707_p1 = $signed(arg_V_read_assign_3_fu_11694_p4);

assign sext_ln700_10_fu_11897_p1 = mul_ln1352_15_fu_11891_p2;

assign sext_ln700_11_fu_12104_p1 = $signed(add_ln700_14_reg_17807);

assign sext_ln700_1_fu_11717_p1 = mul_ln1352_3_fu_11711_p2;

assign sext_ln700_2_fu_12050_p1 = $signed(add_ln700_2_reg_17777);

assign sext_ln700_3_fu_12059_p1 = mul_ln1352_5_reg_17782;

assign sext_ln700_4_fu_11777_p1 = mul_ln1352_7_fu_11771_p2;

assign sext_ln700_5_fu_12068_p1 = $signed(add_ln700_6_reg_17787);

assign sext_ln700_6_fu_12077_p1 = mul_ln1352_9_reg_17792;

assign sext_ln700_7_fu_11837_p1 = mul_ln1352_11_fu_11831_p2;

assign sext_ln700_8_fu_12086_p1 = $signed(add_ln700_10_reg_17797);

assign sext_ln700_9_fu_12095_p1 = mul_ln1352_13_reg_17802;

assign sext_ln700_fu_12041_p1 = mul_ln1352_1_reg_17772;

assign sf_fu_11606_p2 = (32'd1 + sf_1_fu_1406);

assign threshs_m_thresholds_10_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_11_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_12_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_13_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_14_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_15_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_16_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_17_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_18_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_19_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_1_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_20_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_21_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_22_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_23_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_24_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_25_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_26_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_27_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_28_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_29_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_2_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_30_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_31_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_32_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_33_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_34_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_35_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_36_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_37_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_38_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_39_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_3_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_40_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_41_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_42_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_43_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_44_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_45_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_46_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_47_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_48_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_49_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_4_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_50_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_51_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_52_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_53_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_54_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_55_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_5_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_6_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_7_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_8_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_9_address0 = zext_ln142_fu_11916_p1;

assign threshs_m_thresholds_address0 = zext_ln142_fu_11916_p1;

assign trunc_ln321_fu_8559_p1 = sf_1_fu_1406[9:0];

assign trunc_ln647_1_fu_11623_p1 = ap_phi_reg_pp0_iter1_act_m_val_V_reg_4476[3:0];

assign trunc_ln647_fu_11452_p1 = weight_V_V_TDATA[3:0];

assign xor_ln899_10_fu_12715_p2 = (icmp_ln899_10_reg_18142 ^ 1'd1);

assign xor_ln899_11_fu_12724_p2 = (icmp_ln899_11_reg_18147 ^ 1'd1);

assign xor_ln899_12_fu_12733_p2 = (icmp_ln899_12_reg_18152 ^ 1'd1);

assign xor_ln899_13_fu_12742_p2 = (icmp_ln899_13_reg_18157 ^ 1'd1);

assign xor_ln899_14_fu_12861_p2 = (icmp_ln899_14_reg_18162 ^ 1'd1);

assign xor_ln899_15_fu_12870_p2 = (icmp_ln899_15_reg_18167 ^ 1'd1);

assign xor_ln899_16_fu_12879_p2 = (icmp_ln899_16_reg_18172 ^ 1'd1);

assign xor_ln899_17_fu_12888_p2 = (icmp_ln899_17_reg_18177 ^ 1'd1);

assign xor_ln899_18_fu_12897_p2 = (icmp_ln899_18_reg_18182 ^ 1'd1);

assign xor_ln899_19_fu_12906_p2 = (icmp_ln899_19_reg_18187 ^ 1'd1);

assign xor_ln899_1_fu_12634_p2 = (icmp_ln899_1_reg_18097 ^ 1'd1);

assign xor_ln899_20_fu_12915_p2 = (icmp_ln899_20_reg_18192 ^ 1'd1);

assign xor_ln899_21_fu_12924_p2 = (icmp_ln899_21_reg_18197 ^ 1'd1);

assign xor_ln899_22_fu_12933_p2 = (icmp_ln899_22_reg_18202 ^ 1'd1);

assign xor_ln899_23_fu_12942_p2 = (icmp_ln899_23_reg_18207 ^ 1'd1);

assign xor_ln899_24_fu_12951_p2 = (icmp_ln899_24_reg_18212 ^ 1'd1);

assign xor_ln899_25_fu_12960_p2 = (icmp_ln899_25_reg_18217 ^ 1'd1);

assign xor_ln899_26_fu_12969_p2 = (icmp_ln899_26_reg_18222 ^ 1'd1);

assign xor_ln899_27_fu_12978_p2 = (icmp_ln899_27_reg_18227 ^ 1'd1);

assign xor_ln899_28_fu_13097_p2 = (icmp_ln899_28_reg_18232 ^ 1'd1);

assign xor_ln899_29_fu_13106_p2 = (icmp_ln899_29_reg_18237 ^ 1'd1);

assign xor_ln899_2_fu_12643_p2 = (icmp_ln899_2_reg_18102 ^ 1'd1);

assign xor_ln899_30_fu_13115_p2 = (icmp_ln899_30_reg_18242 ^ 1'd1);

assign xor_ln899_31_fu_13124_p2 = (icmp_ln899_31_reg_18247 ^ 1'd1);

assign xor_ln899_32_fu_13133_p2 = (icmp_ln899_32_reg_18252 ^ 1'd1);

assign xor_ln899_33_fu_13142_p2 = (icmp_ln899_33_reg_18257 ^ 1'd1);

assign xor_ln899_34_fu_13151_p2 = (icmp_ln899_34_reg_18262 ^ 1'd1);

assign xor_ln899_35_fu_13160_p2 = (icmp_ln899_35_reg_18267 ^ 1'd1);

assign xor_ln899_36_fu_13169_p2 = (icmp_ln899_36_reg_18272 ^ 1'd1);

assign xor_ln899_37_fu_13178_p2 = (icmp_ln899_37_reg_18277 ^ 1'd1);

assign xor_ln899_38_fu_13187_p2 = (icmp_ln899_38_reg_18282 ^ 1'd1);

assign xor_ln899_39_fu_13196_p2 = (icmp_ln899_39_reg_18287 ^ 1'd1);

assign xor_ln899_3_fu_12652_p2 = (icmp_ln899_3_reg_18107 ^ 1'd1);

assign xor_ln899_40_fu_13205_p2 = (icmp_ln899_40_reg_18292 ^ 1'd1);

assign xor_ln899_41_fu_13214_p2 = (icmp_ln899_41_reg_18297 ^ 1'd1);

assign xor_ln899_42_fu_13333_p2 = (icmp_ln899_42_reg_18302 ^ 1'd1);

assign xor_ln899_43_fu_13342_p2 = (icmp_ln899_43_reg_18307 ^ 1'd1);

assign xor_ln899_44_fu_13351_p2 = (icmp_ln899_44_reg_18312 ^ 1'd1);

assign xor_ln899_45_fu_13360_p2 = (icmp_ln899_45_reg_18317 ^ 1'd1);

assign xor_ln899_46_fu_13369_p2 = (icmp_ln899_46_reg_18322 ^ 1'd1);

assign xor_ln899_47_fu_13378_p2 = (icmp_ln899_47_reg_18327 ^ 1'd1);

assign xor_ln899_48_fu_13387_p2 = (icmp_ln899_48_reg_18332 ^ 1'd1);

assign xor_ln899_49_fu_13396_p2 = (icmp_ln899_49_reg_18337 ^ 1'd1);

assign xor_ln899_4_fu_12661_p2 = (icmp_ln899_4_reg_18112 ^ 1'd1);

assign xor_ln899_50_fu_13405_p2 = (icmp_ln899_50_reg_18342 ^ 1'd1);

assign xor_ln899_51_fu_13414_p2 = (icmp_ln899_51_reg_18347 ^ 1'd1);

assign xor_ln899_52_fu_13423_p2 = (icmp_ln899_52_reg_18352 ^ 1'd1);

assign xor_ln899_53_fu_13432_p2 = (icmp_ln899_53_reg_18357 ^ 1'd1);

assign xor_ln899_54_fu_13441_p2 = (icmp_ln899_54_reg_18362 ^ 1'd1);

assign xor_ln899_55_fu_13450_p2 = (icmp_ln899_55_reg_18367 ^ 1'd1);

assign xor_ln899_5_fu_12670_p2 = (icmp_ln899_5_reg_18117 ^ 1'd1);

assign xor_ln899_6_fu_12679_p2 = (icmp_ln899_6_reg_18122 ^ 1'd1);

assign xor_ln899_7_fu_12688_p2 = (icmp_ln899_7_reg_18127 ^ 1'd1);

assign xor_ln899_8_fu_12697_p2 = (icmp_ln899_8_reg_18132 ^ 1'd1);

assign xor_ln899_9_fu_12706_p2 = (icmp_ln899_9_reg_18137 ^ 1'd1);

assign xor_ln899_fu_12625_p2 = (icmp_ln899_reg_18092 ^ 1'd1);

assign zext_ln142_10_fu_12711_p1 = xor_ln899_9_fu_12706_p2;

assign zext_ln142_11_fu_12720_p1 = xor_ln899_10_fu_12715_p2;

assign zext_ln142_12_fu_12729_p1 = xor_ln899_11_fu_12724_p2;

assign zext_ln142_13_fu_12738_p1 = xor_ln899_12_fu_12733_p2;

assign zext_ln142_14_fu_12866_p1 = xor_ln899_14_fu_12861_p2;

assign zext_ln142_15_fu_12875_p1 = xor_ln899_15_fu_12870_p2;

assign zext_ln142_16_fu_12884_p1 = xor_ln899_16_fu_12879_p2;

assign zext_ln142_17_fu_12893_p1 = xor_ln899_17_fu_12888_p2;

assign zext_ln142_18_fu_12902_p1 = xor_ln899_18_fu_12897_p2;

assign zext_ln142_19_fu_12911_p1 = xor_ln899_19_fu_12906_p2;

assign zext_ln142_1_fu_12630_p1 = xor_ln899_fu_12625_p2;

assign zext_ln142_20_fu_12920_p1 = xor_ln899_20_fu_12915_p2;

assign zext_ln142_21_fu_12929_p1 = xor_ln899_21_fu_12924_p2;

assign zext_ln142_22_fu_12938_p1 = xor_ln899_22_fu_12933_p2;

assign zext_ln142_23_fu_12947_p1 = xor_ln899_23_fu_12942_p2;

assign zext_ln142_24_fu_12956_p1 = xor_ln899_24_fu_12951_p2;

assign zext_ln142_25_fu_12965_p1 = xor_ln899_25_fu_12960_p2;

assign zext_ln142_26_fu_12974_p1 = xor_ln899_26_fu_12969_p2;

assign zext_ln142_27_fu_13102_p1 = xor_ln899_28_fu_13097_p2;

assign zext_ln142_28_fu_13111_p1 = xor_ln899_29_fu_13106_p2;

assign zext_ln142_29_fu_13120_p1 = xor_ln899_30_fu_13115_p2;

assign zext_ln142_2_fu_12639_p1 = xor_ln899_1_fu_12634_p2;

assign zext_ln142_30_fu_13129_p1 = xor_ln899_31_fu_13124_p2;

assign zext_ln142_31_fu_13138_p1 = xor_ln899_32_fu_13133_p2;

assign zext_ln142_32_fu_13147_p1 = xor_ln899_33_fu_13142_p2;

assign zext_ln142_33_fu_13156_p1 = xor_ln899_34_fu_13151_p2;

assign zext_ln142_34_fu_13165_p1 = xor_ln899_35_fu_13160_p2;

assign zext_ln142_35_fu_13174_p1 = xor_ln899_36_fu_13169_p2;

assign zext_ln142_36_fu_13183_p1 = xor_ln899_37_fu_13178_p2;

assign zext_ln142_37_fu_13192_p1 = xor_ln899_38_fu_13187_p2;

assign zext_ln142_38_fu_13201_p1 = xor_ln899_39_fu_13196_p2;

assign zext_ln142_39_fu_13210_p1 = xor_ln899_40_fu_13205_p2;

assign zext_ln142_3_fu_12648_p1 = xor_ln899_2_fu_12643_p2;

assign zext_ln142_40_fu_13338_p1 = xor_ln899_42_fu_13333_p2;

assign zext_ln142_41_fu_13347_p1 = xor_ln899_43_fu_13342_p2;

assign zext_ln142_42_fu_13356_p1 = xor_ln899_44_fu_13351_p2;

assign zext_ln142_43_fu_13365_p1 = xor_ln899_45_fu_13360_p2;

assign zext_ln142_44_fu_13374_p1 = xor_ln899_46_fu_13369_p2;

assign zext_ln142_45_fu_13383_p1 = xor_ln899_47_fu_13378_p2;

assign zext_ln142_46_fu_13392_p1 = xor_ln899_48_fu_13387_p2;

assign zext_ln142_47_fu_13401_p1 = xor_ln899_49_fu_13396_p2;

assign zext_ln142_48_fu_13410_p1 = xor_ln899_50_fu_13405_p2;

assign zext_ln142_49_fu_13419_p1 = xor_ln899_51_fu_13414_p2;

assign zext_ln142_4_fu_12657_p1 = xor_ln899_3_fu_12652_p2;

assign zext_ln142_50_fu_13428_p1 = xor_ln899_52_fu_13423_p2;

assign zext_ln142_51_fu_13437_p1 = xor_ln899_53_fu_13432_p2;

assign zext_ln142_52_fu_13446_p1 = xor_ln899_54_fu_13441_p2;

assign zext_ln142_5_fu_12666_p1 = xor_ln899_4_fu_12661_p2;

assign zext_ln142_6_fu_12675_p1 = xor_ln899_5_fu_12670_p2;

assign zext_ln142_7_fu_12684_p1 = xor_ln899_6_fu_12679_p2;

assign zext_ln142_8_fu_12693_p1 = xor_ln899_7_fu_12688_p2;

assign zext_ln142_9_fu_12702_p1 = xor_ln899_8_fu_12697_p2;

assign zext_ln142_fu_11916_p1 = nf_assign_fu_3714;

assign zext_ln700_10_fu_12999_p1 = add_ln700_30_fu_12993_p2;

assign zext_ln700_11_fu_13009_p1 = add_ln700_31_fu_13003_p2;

assign zext_ln700_12_fu_13019_p1 = add_ln700_32_fu_13013_p2;

assign zext_ln700_13_fu_13035_p1 = add_ln700_34_fu_13029_p2;

assign zext_ln700_14_fu_13051_p1 = add_ln700_36_fu_13045_p2;

assign zext_ln700_15_fu_13061_p1 = add_ln700_37_fu_13055_p2;

assign zext_ln700_16_fu_13071_p1 = add_ln700_38_fu_13065_p2;

assign zext_ln700_17_fu_13087_p1 = add_ln700_40_fu_13081_p2;

assign zext_ln700_18_fu_13219_p1 = xor_ln899_41_fu_13214_p2;

assign zext_ln700_19_fu_13235_p1 = add_ln700_43_fu_13229_p2;

assign zext_ln700_1_fu_12763_p1 = add_ln700_17_fu_12757_p2;

assign zext_ln700_20_fu_13245_p1 = add_ln700_44_fu_13239_p2;

assign zext_ln700_21_fu_13255_p1 = add_ln700_45_fu_13249_p2;

assign zext_ln700_22_fu_13271_p1 = add_ln700_47_fu_13265_p2;

assign zext_ln700_23_fu_13287_p1 = add_ln700_49_fu_13281_p2;

assign zext_ln700_24_fu_13297_p1 = add_ln700_50_fu_13291_p2;

assign zext_ln700_25_fu_13307_p1 = add_ln700_51_fu_13301_p2;

assign zext_ln700_26_fu_13323_p1 = add_ln700_53_fu_13317_p2;

assign zext_ln700_27_fu_13455_p1 = xor_ln899_55_fu_13450_p2;

assign zext_ln700_28_fu_13471_p1 = add_ln700_56_fu_13465_p2;

assign zext_ln700_29_fu_13481_p1 = add_ln700_57_fu_13475_p2;

assign zext_ln700_2_fu_12773_p1 = add_ln700_18_fu_12767_p2;

assign zext_ln700_30_fu_13491_p1 = add_ln700_58_fu_13485_p2;

assign zext_ln700_31_fu_13507_p1 = add_ln700_60_fu_13501_p2;

assign zext_ln700_32_fu_13523_p1 = add_ln700_62_fu_13517_p2;

assign zext_ln700_33_fu_13533_p1 = add_ln700_63_fu_13527_p2;

assign zext_ln700_34_fu_13543_p1 = add_ln700_64_fu_13537_p2;

assign zext_ln700_35_fu_13559_p1 = add_ln700_66_fu_13553_p2;

assign zext_ln700_3_fu_12783_p1 = add_ln700_19_fu_12777_p2;

assign zext_ln700_4_fu_12799_p1 = add_ln700_21_fu_12793_p2;

assign zext_ln700_5_fu_12815_p1 = add_ln700_23_fu_12809_p2;

assign zext_ln700_6_fu_12825_p1 = add_ln700_24_fu_12819_p2;

assign zext_ln700_7_fu_12835_p1 = add_ln700_25_fu_12829_p2;

assign zext_ln700_8_fu_12851_p1 = add_ln700_27_fu_12845_p2;

assign zext_ln700_9_fu_12983_p1 = xor_ln899_27_fu_12978_p2;

assign zext_ln700_fu_12747_p1 = xor_ln899_13_fu_12742_p2;

endmodule //StreamingFCLayer_Batch_1_Matrix_Vector_Activa
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Act3i2.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Act3i2_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Act3i2_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Act3i2(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Act3i2_rom StreamingFCLayer_Batch_3_Matrix_Vector_Act3i2_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_BatckbM.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_BatckbM_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_BatckbM_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_BatckbM(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_BatckbM_rom Thresholding_Batch_2_Thresholding_BatckbM_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc1C.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcc1C_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc1C_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcc1C(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcc1C_rom Thresholding_Batch_0_Thresholding_Batcc1C_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc2C.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcc2C_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcc2C_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcc2C(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcc2C_rom Thresholding_Batch_0_Thresholding_Batcc2C_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/7fe4/hdl/verilog/StreamingDataWidthConverter_Batch_3_StreamingDataWidthConverter_Batch_3.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingDataWidthConverter_Batch_3_StreamingDataWidthConverter_Batch_3,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=5.025000,HLS_SYN_LAT=133,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=116,HLS_SYN_LUT=225,HLS_VERSION=2020_1_1}" *)

module StreamingDataWidthConverter_Batch_3_StreamingDataWidthConverter_Batch_3 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_start;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_done;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_idle;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_ready;
wire    grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
wire   [31:0] grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY;
reg    grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [15:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_StreamingDataWidthCo_1_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingDataWidthConverter_Batch_3_StreamingDataWidthCo_1 grp_StreamingDataWidthCo_1_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_StreamingDataWidthCo_1_fu_26_ap_start),
    .ap_done(grp_StreamingDataWidthCo_1_fu_26_ap_done),
    .ap_idle(grp_StreamingDataWidthCo_1_fu_26_ap_idle),
    .ap_ready(grp_StreamingDataWidthCo_1_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 32 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .vld_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_StreamingDataWidthCo_1_fu_26_ap_ready == 1'b1)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_StreamingDataWidthCo_1_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_StreamingDataWidthCo_1_fu_26_ap_start = grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;

assign grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingDataWidthConverter_Batch_3_StreamingDataWidthConverter_Batch_3
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/46bc/StreamingFIFO_19.v


module StreamingFIFO_19(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [7:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(8)
)
StreamingFIFO_19_StreamingFIFO_19
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/a3f1/hdl/verilog/ConvolutionInputGenerator_1_ConvolutionInputGenerator_1.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="ConvolutionInputGenerator_1_ConvolutionInputGenerator_1,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=7.832750,HLS_SYN_LAT=1157,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=473,HLS_SYN_LUT=1561,HLS_VERSION=2020_1_1}" *)

module ConvolutionInputGenerator_1_ConvolutionInputGenerator_1 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_ConvolutionInputGene_1_fu_26_ap_start;
wire    grp_ConvolutionInputGene_1_fu_26_ap_done;
wire    grp_ConvolutionInputGene_1_fu_26_ap_idle;
wire    grp_ConvolutionInputGene_1_fu_26_ap_ready;
wire    grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY;
wire   [15:0] grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA;
wire    grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID;
wire    grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY;
reg    grp_ConvolutionInputGene_1_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [15:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_ConvolutionInputGene_1_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

ConvolutionInputGenerator_1_ConvolutionInputGene_1 grp_ConvolutionInputGene_1_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_ConvolutionInputGene_1_fu_26_ap_start),
    .ap_done(grp_ConvolutionInputGene_1_fu_26_ap_done),
    .ap_idle(grp_ConvolutionInputGene_1_fu_26_ap_idle),
    .ap_ready(grp_ConvolutionInputGene_1_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_ConvolutionInputGene_1_fu_26_out_V_V_TDATA),
    .vld_in(grp_ConvolutionInputGene_1_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_ConvolutionInputGene_1_fu_26_ap_ready == 1'b1)) begin
            grp_ConvolutionInputGene_1_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_ConvolutionInputGene_1_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_ConvolutionInputGene_1_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_ConvolutionInputGene_1_fu_26_ap_start = grp_ConvolutionInputGene_1_fu_26_ap_start_reg;

assign grp_ConvolutionInputGene_1_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //ConvolutionInputGenerator_1_ConvolutionInputGenerator_1
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actzec.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actzec_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_Actzec_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_Actzec(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_Actzec_rom StreamingFCLayer_Batch_1_Matrix_Vector_Actzec_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatceOg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatceOg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 3;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatceOg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatceOg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd3;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatceOg_rom Thresholding_Batch_0_Thresholding_BatceOg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActLf8.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActLf8_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActLf8_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActLf8(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActLf8_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActLf8_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_Thresholding_Batch_1_0/synth/finn_design_Thresholding_Batch_1_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:Thresholding_Batch_1:1.0
// IP Revision: 2101301317

(* X_CORE_INFO = "Thresholding_Batch_1_Thresholding_Batch_1,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_Thresholding_Batch_1_0,Thresholding_Batch_1_Thresholding_Batch_1,{}" *)
(* CORE_GENERATION_INFO = "finn_design_Thresholding_Batch_1_0,Thresholding_Batch_1_Thresholding_Batch_1,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=Thresholding_Batch_1,x_ipVersion=1.0,x_ipCoreRevision=2101301317,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* IP_DEFINITION_SOURCE = "HLS" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_Thresholding_Batch_1_0 (
  ap_clk,
  ap_rst_n,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  in0_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY,
  out_V_V_TDATA
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, ASSOCIATED_RESET ap_rst_n, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 3, TUSER_WIDTH 0, LAYERED_METADATA undef, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [23 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TUSER_WIDTH 0, TDEST_WIDTH 0, TID_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;

  Thresholding_Batch_1_Thresholding_Batch_1 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcxdS.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcxdS_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 5;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcxdS_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcxdS(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd5;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcxdS_rom Thresholding_Batch_0_Thresholding_BatcxdS_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActHfu.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActHfu_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActHfu_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActHfu(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActHfu_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActHfu_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8ee6/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbek.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbek_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbek_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbek(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbek_rom Thresholding_Batch_0_Thresholding_Batcbek_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccXB.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccXB_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccXB_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccXB(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccXB_rom Thresholding_Batch_0_Thresholding_BatccXB_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actvdy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actvdy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 15;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Actvdy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Actvdy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd15;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Actvdy_rom StreamingFCLayer_Batch_3_Matrix_Vector_Actvdy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccwx.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batccwx_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batccwx_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batccwx(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batccwx_rom Thresholding_Batch_0_Thresholding_Batccwx_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActNgs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActNgs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActNgs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActNgs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActNgs_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActNgs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActUhA.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActUhA_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActUhA_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActUhA(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActUhA_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActUhA_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcvdy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcvdy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 5;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcvdy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcvdy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd5;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcvdy_rom Thresholding_Batch_0_Thresholding_Batcvdy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ip/finn_design_StreamingFIFO_1_0/synth/finn_design_StreamingFIFO_1_0.v

// (c) Copyright 1995-2021 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// 
// DO NOT MODIFY THIS FILE.


// IP VLNV: xilinx.com:hls:StreamingFIFO_1:1.0
// IP Revision: 2

(* X_CORE_INFO = "StreamingFIFO_1,Vivado 2020.1.1" *)
(* CHECK_LICENSE_TYPE = "finn_design_StreamingFIFO_1_0,StreamingFIFO_1,{}" *)
(* CORE_GENERATION_INFO = "finn_design_StreamingFIFO_1_0,StreamingFIFO_1,{x_ipProduct=Vivado 2020.1.1,x_ipVendor=xilinx.com,x_ipLibrary=hls,x_ipName=StreamingFIFO_1,x_ipVersion=1.0,x_ipCoreRevision=2,x_ipLanguage=VERILOG,x_ipSimLanguage=MIXED}" *)
(* DowngradeIPIdentifiedWarnings = "yes" *)
module finn_design_StreamingFIFO_1_0 (
  ap_clk,
  ap_rst_n,
  count,
  in0_V_V_TDATA,
  in0_V_V_TVALID,
  in0_V_V_TREADY,
  out_V_V_TDATA,
  out_V_V_TVALID,
  out_V_V_TREADY
);

(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_clk, ASSOCIATED_BUSIF in0_V_V:out_V_V, FREQ_HZ 100000000.000000, FREQ_TOLERANCE_HZ 0, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ap_clk CLK" *)
input wire ap_clk;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME ap_rst_n, POLARITY ACTIVE_LOW, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 ap_rst_n RST" *)
input wire ap_rst_n;
output wire [13 : 0] count;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TDATA" *)
input wire [7 : 0] in0_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TVALID" *)
input wire in0_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME in0_V_V, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 in0_V_V TREADY" *)
output wire in0_V_V_TREADY;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TDATA" *)
output wire [7 : 0] out_V_V_TDATA;
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TVALID" *)
output wire out_V_V_TVALID;
(* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME out_V_V, TDATA_NUM_BYTES 1, TDEST_WIDTH 0, TID_WIDTH 0, TUSER_WIDTH 0, HAS_TREADY 1, HAS_TSTRB 0, HAS_TKEEP 0, HAS_TLAST 0, FREQ_HZ 100000000.000000, PHASE 0.000, CLK_DOMAIN finn_design_ap_clk_0, LAYERED_METADATA undef, INSERT_VIP 0" *)
(* X_INTERFACE_INFO = "xilinx.com:interface:axis:1.0 out_V_V TREADY" *)
input wire out_V_V_TREADY;

  StreamingFIFO_1 inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .count(count),
    .in0_V_V_TDATA(in0_V_V_TDATA),
    .in0_V_V_TVALID(in0_V_V_TVALID),
    .in0_V_V_TREADY(in0_V_V_TREADY),
    .out_V_V_TDATA(out_V_V_TDATA),
    .out_V_V_TVALID(out_V_V_TVALID),
    .out_V_V_TREADY(out_V_V_TREADY)
  );
endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActShg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActShg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActShg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActShg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActShg_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActShg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActFfa.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActFfa_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActFfa_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActFfa(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActFfa_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActFfa_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbck.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbck_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbck_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbck(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbck_rom Thresholding_Batch_0_Thresholding_Batcbck_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_StreamingFCLayer_5jm.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module StreamingFCLayer_Batch_4_StreamingFCLayer_5jm #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH       = 32,
    din5_WIDTH       = 32,
    din6_WIDTH       = 32,
    din7_WIDTH       = 32,
    din8_WIDTH       = 32,
    din9_WIDTH       = 32,
    din10_WIDTH       = 32,
    din11_WIDTH       = 32,
    din12_WIDTH       = 32,
    din13_WIDTH       = 32,
    din14_WIDTH       = 32,
    din15_WIDTH       = 32,
    din16_WIDTH       = 32,
    din17_WIDTH       = 32,
    din18_WIDTH       = 32,
    din19_WIDTH       = 32,
    din20_WIDTH       = 32,
    din21_WIDTH       = 32,
    din22_WIDTH       = 32,
    din23_WIDTH       = 32,
    din24_WIDTH       = 32,
    din25_WIDTH       = 32,
    din26_WIDTH       = 32,
    din27_WIDTH       = 32,
    din28_WIDTH       = 32,
    din29_WIDTH       = 32,
    din30_WIDTH       = 32,
    din31_WIDTH       = 32,
    din32_WIDTH       = 32,
    din33_WIDTH       = 32,
    din34_WIDTH       = 32,
    din35_WIDTH       = 32,
    din36_WIDTH       = 32,
    din37_WIDTH       = 32,
    din38_WIDTH       = 32,
    din39_WIDTH       = 32,
    din40_WIDTH       = 32,
    din41_WIDTH       = 32,
    din42_WIDTH       = 32,
    din43_WIDTH       = 32,
    din44_WIDTH       = 32,
    din45_WIDTH       = 32,
    din46_WIDTH       = 32,
    din47_WIDTH       = 32,
    din48_WIDTH       = 32,
    din49_WIDTH       = 32,
    din50_WIDTH       = 32,
    din51_WIDTH       = 32,
    din52_WIDTH       = 32,
    din53_WIDTH       = 32,
    din54_WIDTH       = 32,
    din55_WIDTH       = 32,
    din56_WIDTH       = 32,
    din57_WIDTH       = 32,
    din58_WIDTH       = 32,
    din59_WIDTH       = 32,
    din60_WIDTH       = 32,
    din61_WIDTH       = 32,
    din62_WIDTH       = 32,
    din63_WIDTH       = 32,
    din64_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [31 : 0]     din0,
    input  [31 : 0]     din1,
    input  [31 : 0]     din2,
    input  [31 : 0]     din3,
    input  [31 : 0]     din4,
    input  [31 : 0]     din5,
    input  [31 : 0]     din6,
    input  [31 : 0]     din7,
    input  [31 : 0]     din8,
    input  [31 : 0]     din9,
    input  [31 : 0]     din10,
    input  [31 : 0]     din11,
    input  [31 : 0]     din12,
    input  [31 : 0]     din13,
    input  [31 : 0]     din14,
    input  [31 : 0]     din15,
    input  [31 : 0]     din16,
    input  [31 : 0]     din17,
    input  [31 : 0]     din18,
    input  [31 : 0]     din19,
    input  [31 : 0]     din20,
    input  [31 : 0]     din21,
    input  [31 : 0]     din22,
    input  [31 : 0]     din23,
    input  [31 : 0]     din24,
    input  [31 : 0]     din25,
    input  [31 : 0]     din26,
    input  [31 : 0]     din27,
    input  [31 : 0]     din28,
    input  [31 : 0]     din29,
    input  [31 : 0]     din30,
    input  [31 : 0]     din31,
    input  [31 : 0]     din32,
    input  [31 : 0]     din33,
    input  [31 : 0]     din34,
    input  [31 : 0]     din35,
    input  [31 : 0]     din36,
    input  [31 : 0]     din37,
    input  [31 : 0]     din38,
    input  [31 : 0]     din39,
    input  [31 : 0]     din40,
    input  [31 : 0]     din41,
    input  [31 : 0]     din42,
    input  [31 : 0]     din43,
    input  [31 : 0]     din44,
    input  [31 : 0]     din45,
    input  [31 : 0]     din46,
    input  [31 : 0]     din47,
    input  [31 : 0]     din48,
    input  [31 : 0]     din49,
    input  [31 : 0]     din50,
    input  [31 : 0]     din51,
    input  [31 : 0]     din52,
    input  [31 : 0]     din53,
    input  [31 : 0]     din54,
    input  [31 : 0]     din55,
    input  [31 : 0]     din56,
    input  [31 : 0]     din57,
    input  [31 : 0]     din58,
    input  [31 : 0]     din59,
    input  [31 : 0]     din60,
    input  [31 : 0]     din61,
    input  [31 : 0]     din62,
    input  [31 : 0]     din63,
    input  [5 : 0]    din64,
    output [31 : 0]   dout);

// puts internal signals
wire [5 : 0]     sel;
// level 1 signals
wire [31 : 0]         mux_1_0;
wire [31 : 0]         mux_1_1;
wire [31 : 0]         mux_1_2;
wire [31 : 0]         mux_1_3;
wire [31 : 0]         mux_1_4;
wire [31 : 0]         mux_1_5;
wire [31 : 0]         mux_1_6;
wire [31 : 0]         mux_1_7;
wire [31 : 0]         mux_1_8;
wire [31 : 0]         mux_1_9;
wire [31 : 0]         mux_1_10;
wire [31 : 0]         mux_1_11;
wire [31 : 0]         mux_1_12;
wire [31 : 0]         mux_1_13;
wire [31 : 0]         mux_1_14;
wire [31 : 0]         mux_1_15;
wire [31 : 0]         mux_1_16;
wire [31 : 0]         mux_1_17;
wire [31 : 0]         mux_1_18;
wire [31 : 0]         mux_1_19;
wire [31 : 0]         mux_1_20;
wire [31 : 0]         mux_1_21;
wire [31 : 0]         mux_1_22;
wire [31 : 0]         mux_1_23;
wire [31 : 0]         mux_1_24;
wire [31 : 0]         mux_1_25;
wire [31 : 0]         mux_1_26;
wire [31 : 0]         mux_1_27;
wire [31 : 0]         mux_1_28;
wire [31 : 0]         mux_1_29;
wire [31 : 0]         mux_1_30;
wire [31 : 0]         mux_1_31;
// level 2 signals
wire [31 : 0]         mux_2_0;
wire [31 : 0]         mux_2_1;
wire [31 : 0]         mux_2_2;
wire [31 : 0]         mux_2_3;
wire [31 : 0]         mux_2_4;
wire [31 : 0]         mux_2_5;
wire [31 : 0]         mux_2_6;
wire [31 : 0]         mux_2_7;
wire [31 : 0]         mux_2_8;
wire [31 : 0]         mux_2_9;
wire [31 : 0]         mux_2_10;
wire [31 : 0]         mux_2_11;
wire [31 : 0]         mux_2_12;
wire [31 : 0]         mux_2_13;
wire [31 : 0]         mux_2_14;
wire [31 : 0]         mux_2_15;
// level 3 signals
wire [31 : 0]         mux_3_0;
wire [31 : 0]         mux_3_1;
wire [31 : 0]         mux_3_2;
wire [31 : 0]         mux_3_3;
wire [31 : 0]         mux_3_4;
wire [31 : 0]         mux_3_5;
wire [31 : 0]         mux_3_6;
wire [31 : 0]         mux_3_7;
// level 4 signals
wire [31 : 0]         mux_4_0;
wire [31 : 0]         mux_4_1;
wire [31 : 0]         mux_4_2;
wire [31 : 0]         mux_4_3;
// level 5 signals
wire [31 : 0]         mux_5_0;
wire [31 : 0]         mux_5_1;
// level 6 signals
wire [31 : 0]         mux_6_0;

assign sel = din64;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;
assign mux_1_2 = (sel[0] == 0)? din4 : din5;
assign mux_1_3 = (sel[0] == 0)? din6 : din7;
assign mux_1_4 = (sel[0] == 0)? din8 : din9;
assign mux_1_5 = (sel[0] == 0)? din10 : din11;
assign mux_1_6 = (sel[0] == 0)? din12 : din13;
assign mux_1_7 = (sel[0] == 0)? din14 : din15;
assign mux_1_8 = (sel[0] == 0)? din16 : din17;
assign mux_1_9 = (sel[0] == 0)? din18 : din19;
assign mux_1_10 = (sel[0] == 0)? din20 : din21;
assign mux_1_11 = (sel[0] == 0)? din22 : din23;
assign mux_1_12 = (sel[0] == 0)? din24 : din25;
assign mux_1_13 = (sel[0] == 0)? din26 : din27;
assign mux_1_14 = (sel[0] == 0)? din28 : din29;
assign mux_1_15 = (sel[0] == 0)? din30 : din31;
assign mux_1_16 = (sel[0] == 0)? din32 : din33;
assign mux_1_17 = (sel[0] == 0)? din34 : din35;
assign mux_1_18 = (sel[0] == 0)? din36 : din37;
assign mux_1_19 = (sel[0] == 0)? din38 : din39;
assign mux_1_20 = (sel[0] == 0)? din40 : din41;
assign mux_1_21 = (sel[0] == 0)? din42 : din43;
assign mux_1_22 = (sel[0] == 0)? din44 : din45;
assign mux_1_23 = (sel[0] == 0)? din46 : din47;
assign mux_1_24 = (sel[0] == 0)? din48 : din49;
assign mux_1_25 = (sel[0] == 0)? din50 : din51;
assign mux_1_26 = (sel[0] == 0)? din52 : din53;
assign mux_1_27 = (sel[0] == 0)? din54 : din55;
assign mux_1_28 = (sel[0] == 0)? din56 : din57;
assign mux_1_29 = (sel[0] == 0)? din58 : din59;
assign mux_1_30 = (sel[0] == 0)? din60 : din61;
assign mux_1_31 = (sel[0] == 0)? din62 : din63;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;
assign mux_2_1 = (sel[1] == 0)? mux_1_2 : mux_1_3;
assign mux_2_2 = (sel[1] == 0)? mux_1_4 : mux_1_5;
assign mux_2_3 = (sel[1] == 0)? mux_1_6 : mux_1_7;
assign mux_2_4 = (sel[1] == 0)? mux_1_8 : mux_1_9;
assign mux_2_5 = (sel[1] == 0)? mux_1_10 : mux_1_11;
assign mux_2_6 = (sel[1] == 0)? mux_1_12 : mux_1_13;
assign mux_2_7 = (sel[1] == 0)? mux_1_14 : mux_1_15;
assign mux_2_8 = (sel[1] == 0)? mux_1_16 : mux_1_17;
assign mux_2_9 = (sel[1] == 0)? mux_1_18 : mux_1_19;
assign mux_2_10 = (sel[1] == 0)? mux_1_20 : mux_1_21;
assign mux_2_11 = (sel[1] == 0)? mux_1_22 : mux_1_23;
assign mux_2_12 = (sel[1] == 0)? mux_1_24 : mux_1_25;
assign mux_2_13 = (sel[1] == 0)? mux_1_26 : mux_1_27;
assign mux_2_14 = (sel[1] == 0)? mux_1_28 : mux_1_29;
assign mux_2_15 = (sel[1] == 0)? mux_1_30 : mux_1_31;

// Generate level 3 logic
assign mux_3_0 = (sel[2] == 0)? mux_2_0 : mux_2_1;
assign mux_3_1 = (sel[2] == 0)? mux_2_2 : mux_2_3;
assign mux_3_2 = (sel[2] == 0)? mux_2_4 : mux_2_5;
assign mux_3_3 = (sel[2] == 0)? mux_2_6 : mux_2_7;
assign mux_3_4 = (sel[2] == 0)? mux_2_8 : mux_2_9;
assign mux_3_5 = (sel[2] == 0)? mux_2_10 : mux_2_11;
assign mux_3_6 = (sel[2] == 0)? mux_2_12 : mux_2_13;
assign mux_3_7 = (sel[2] == 0)? mux_2_14 : mux_2_15;

// Generate level 4 logic
assign mux_4_0 = (sel[3] == 0)? mux_3_0 : mux_3_1;
assign mux_4_1 = (sel[3] == 0)? mux_3_2 : mux_3_3;
assign mux_4_2 = (sel[3] == 0)? mux_3_4 : mux_3_5;
assign mux_4_3 = (sel[3] == 0)? mux_3_6 : mux_3_7;

// Generate level 5 logic
assign mux_5_0 = (sel[4] == 0)? mux_4_0 : mux_4_1;
assign mux_5_1 = (sel[4] == 0)? mux_4_2 : mux_4_3;

// Generate level 6 logic
assign mux_6_0 = (sel[5] == 0)? mux_5_0 : mux_5_1;

// output logic
assign dout = mux_6_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/eb12/StreamingFIFO_9.v


module StreamingFIFO_9(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [23:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [23:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(24)
)
StreamingFIFO_9_StreamingFIFO_9
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActWhU.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_ActWhU_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_ActWhU_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_ActWhU(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_ActWhU_rom StreamingFCLayer_Batch_2_Matrix_Vector_ActWhU_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/ca29/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcncg.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_2_Thresholding_Batcncg_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_2_0eb7bn2y/project_Thresholding_Batch_2/sol1/impl/ip/hdl/verilog/Thresholding_Batch_2_Thresholding_Batcncg_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_2_Thresholding_Batcncg(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_2_Thresholding_Batcncg_rom Thresholding_Batch_2_Thresholding_Batcncg_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actsc4.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actsc4_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_Actsc4_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_Actsc4(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_Actsc4_rom StreamingFCLayer_Batch_4_Matrix_Vector_Actsc4_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActEe0.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActEe0_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActEe0_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActEe0(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActEe0_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActEe0_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Act0iy.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Act0iy_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_Act0iy_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_Act0iy(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_Act0iy_rom StreamingFCLayer_Batch_3_Matrix_Vector_Act0iy_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActBew.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActBew_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActBew_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActBew(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActBew_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActBew_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_Batch.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module Thresholding_Batch_1_Thresholding_Batch (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        in_V_V_TDATA,
        in_V_V_TVALID,
        in_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state5 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [23:0] in_V_V_TDATA;
input   in_V_V_TVALID;
output   in_V_V_TREADY;
output  [7:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_V_V_TREADY;
reg out_V_V_TVALID;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [6:0] threshs_m_thresholds_13_address0;
reg    threshs_m_thresholds_13_ce0;
wire   [18:0] threshs_m_thresholds_13_q0;
wire   [6:0] threshs_m_thresholds_12_address0;
reg    threshs_m_thresholds_12_ce0;
wire   [18:0] threshs_m_thresholds_12_q0;
wire   [6:0] threshs_m_thresholds_7_address0;
reg    threshs_m_thresholds_7_ce0;
wire   [18:0] threshs_m_thresholds_7_q0;
wire   [6:0] threshs_m_thresholds_6_address0;
reg    threshs_m_thresholds_6_ce0;
wire   [18:0] threshs_m_thresholds_6_q0;
wire   [6:0] threshs_m_thresholds_5_address0;
reg    threshs_m_thresholds_5_ce0;
wire   [18:0] threshs_m_thresholds_5_q0;
wire   [6:0] threshs_m_thresholds_4_address0;
reg    threshs_m_thresholds_4_ce0;
wire   [18:0] threshs_m_thresholds_4_q0;
wire   [6:0] threshs_m_thresholds_3_address0;
reg    threshs_m_thresholds_3_ce0;
wire   [18:0] threshs_m_thresholds_3_q0;
wire   [6:0] threshs_m_thresholds_2_address0;
reg    threshs_m_thresholds_2_ce0;
wire   [18:0] threshs_m_thresholds_2_q0;
wire   [6:0] threshs_m_thresholds_1_address0;
reg    threshs_m_thresholds_1_ce0;
wire   [18:0] threshs_m_thresholds_1_q0;
wire   [6:0] threshs_m_thresholds_address0;
reg    threshs_m_thresholds_ce0;
wire   [18:0] threshs_m_thresholds_q0;
wire   [6:0] threshs_m_thresholds_11_address0;
reg    threshs_m_thresholds_11_ce0;
wire   [18:0] threshs_m_thresholds_11_q0;
wire   [6:0] threshs_m_thresholds_10_address0;
reg    threshs_m_thresholds_10_ce0;
wire   [18:0] threshs_m_thresholds_10_q0;
wire   [6:0] threshs_m_thresholds_9_address0;
reg    threshs_m_thresholds_9_ce0;
wire   [18:0] threshs_m_thresholds_9_q0;
wire   [6:0] threshs_m_thresholds_8_address0;
reg    threshs_m_thresholds_8_ce0;
wire   [18:0] threshs_m_thresholds_8_q0;
reg    in_V_V_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_pp0_stage0;
wire   [0:0] icmp_ln221_fu_299_p2;
reg    out_V_V_TDATA_blk_n;
reg    ap_enable_reg_pp0_iter2;
reg   [0:0] icmp_ln221_reg_720;
reg   [0:0] icmp_ln221_reg_720_pp0_iter1_reg;
reg   [31:0] nf_assign_reg_277;
reg   [13:0] i_0_reg_288;
reg    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
reg    ap_block_state4_io;
reg    ap_block_pp0_stage0_11001;
wire   [13:0] i_fu_305_p2;
reg   [23:0] tmp_V_1_reg_729;
wire   [31:0] nf_1_fu_341_p3;
wire   [0:0] icmp_ln899_fu_353_p2;
reg   [0:0] icmp_ln899_reg_822;
wire   [0:0] icmp_ln899_1_fu_362_p2;
reg   [0:0] icmp_ln899_1_reg_827;
wire   [0:0] icmp_ln899_2_fu_371_p2;
reg   [0:0] icmp_ln899_2_reg_832;
wire   [0:0] icmp_ln899_3_fu_380_p2;
reg   [0:0] icmp_ln899_3_reg_837;
wire   [0:0] icmp_ln899_4_fu_389_p2;
reg   [0:0] icmp_ln899_4_reg_842;
wire   [0:0] icmp_ln899_5_fu_398_p2;
reg   [0:0] icmp_ln899_5_reg_847;
wire   [0:0] icmp_ln899_6_fu_407_p2;
reg   [0:0] icmp_ln899_6_reg_852;
wire   [0:0] xor_ln899_7_fu_421_p2;
reg   [0:0] xor_ln899_7_reg_857;
wire   [0:0] xor_ln899_8_fu_436_p2;
reg   [0:0] xor_ln899_8_reg_862;
wire   [0:0] xor_ln899_9_fu_451_p2;
reg   [0:0] xor_ln899_9_reg_867;
wire   [0:0] icmp_ln899_10_fu_461_p2;
reg   [0:0] icmp_ln899_10_reg_872;
wire   [0:0] icmp_ln899_11_fu_470_p2;
reg   [0:0] icmp_ln899_11_reg_877;
wire   [0:0] icmp_ln899_12_fu_479_p2;
reg   [0:0] icmp_ln899_12_reg_882;
wire   [0:0] icmp_ln899_13_fu_488_p2;
reg   [0:0] icmp_ln899_13_reg_887;
reg    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
wire   [63:0] zext_ln142_fu_311_p1;
reg    ap_block_pp0_stage0_01001;
wire   [31:0] nf_fu_329_p2;
wire   [0:0] icmp_ln235_fu_335_p2;
wire  signed [23:0] sext_ln142_fu_349_p1;
wire  signed [23:0] sext_ln142_1_fu_358_p1;
wire  signed [23:0] sext_ln142_2_fu_367_p1;
wire  signed [23:0] sext_ln142_3_fu_376_p1;
wire  signed [23:0] sext_ln142_4_fu_385_p1;
wire  signed [23:0] sext_ln142_5_fu_394_p1;
wire  signed [23:0] sext_ln142_6_fu_403_p1;
wire  signed [23:0] sext_ln142_7_fu_412_p1;
wire   [0:0] icmp_ln899_7_fu_416_p2;
wire  signed [23:0] sext_ln142_8_fu_427_p1;
wire   [0:0] icmp_ln899_8_fu_431_p2;
wire  signed [23:0] sext_ln142_9_fu_442_p1;
wire   [0:0] icmp_ln899_9_fu_446_p2;
wire  signed [23:0] sext_ln142_10_fu_457_p1;
wire  signed [23:0] sext_ln142_11_fu_466_p1;
wire  signed [23:0] sext_ln142_12_fu_475_p1;
wire  signed [23:0] sext_ln142_13_fu_484_p1;
wire   [0:0] xor_ln899_fu_493_p2;
wire   [0:0] xor_ln899_1_fu_506_p2;
wire   [0:0] xor_ln899_2_fu_515_p2;
wire   [0:0] xor_ln899_3_fu_524_p2;
wire   [0:0] xor_ln899_4_fu_533_p2;
wire   [0:0] xor_ln899_5_fu_542_p2;
wire   [0:0] xor_ln899_6_fu_551_p2;
wire   [0:0] xor_ln899_10_fu_569_p2;
wire   [0:0] xor_ln899_11_fu_578_p2;
wire   [0:0] xor_ln899_12_fu_587_p2;
wire   [0:0] xor_ln899_13_fu_596_p2;
wire   [1:0] zext_ln142_1_fu_511_p1;
wire   [1:0] zext_ln142_2_fu_520_p1;
wire   [1:0] add_ln700_fu_605_p2;
wire   [3:0] zext_ln700_1_fu_611_p1;
wire   [3:0] select_ln700_fu_498_p3;
wire   [1:0] zext_ln142_3_fu_529_p1;
wire   [1:0] zext_ln142_4_fu_538_p1;
wire   [1:0] add_ln700_2_fu_621_p2;
wire   [1:0] zext_ln142_5_fu_547_p1;
wire   [1:0] zext_ln142_6_fu_556_p1;
wire   [1:0] add_ln700_3_fu_631_p2;
wire   [2:0] zext_ln700_3_fu_637_p1;
wire   [2:0] zext_ln700_2_fu_627_p1;
wire   [2:0] add_ln700_4_fu_641_p2;
wire   [3:0] zext_ln700_4_fu_647_p1;
wire   [3:0] add_ln700_1_fu_615_p2;
wire   [1:0] zext_ln142_8_fu_563_p1;
wire   [1:0] zext_ln142_9_fu_566_p1;
wire   [1:0] add_ln700_6_fu_657_p2;
wire   [1:0] zext_ln142_7_fu_560_p1;
wire   [1:0] add_ln700_7_fu_663_p2;
wire   [1:0] zext_ln142_10_fu_574_p1;
wire   [1:0] zext_ln142_11_fu_583_p1;
wire   [1:0] add_ln700_8_fu_673_p2;
wire   [1:0] zext_ln142_12_fu_592_p1;
wire   [1:0] zext_ln700_fu_601_p1;
wire   [1:0] add_ln700_9_fu_683_p2;
wire   [2:0] zext_ln700_7_fu_689_p1;
wire   [2:0] zext_ln700_6_fu_679_p1;
wire   [2:0] add_ln700_10_fu_693_p2;
wire   [2:0] zext_ln700_5_fu_669_p1;
wire   [2:0] add_ln700_11_fu_699_p2;
wire   [3:0] zext_ln700_8_fu_705_p1;
wire   [3:0] add_ln700_5_fu_651_p2;
wire   [3:0] tmp_V_fu_709_p2;
wire    ap_CS_fsm_state5;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
end

Thresholding_Batch_1_Thresholding_Batcbkb #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_13_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_13_address0),
    .ce0(threshs_m_thresholds_13_ce0),
    .q0(threshs_m_thresholds_13_q0)
);

Thresholding_Batch_1_Thresholding_Batccud #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_12_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_12_address0),
    .ce0(threshs_m_thresholds_12_ce0),
    .q0(threshs_m_thresholds_12_q0)
);

Thresholding_Batch_1_Thresholding_BatcdEe #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_7_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_7_address0),
    .ce0(threshs_m_thresholds_7_ce0),
    .q0(threshs_m_thresholds_7_q0)
);

Thresholding_Batch_1_Thresholding_BatceOg #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_6_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_6_address0),
    .ce0(threshs_m_thresholds_6_ce0),
    .q0(threshs_m_thresholds_6_q0)
);

Thresholding_Batch_1_Thresholding_BatcfYi #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_5_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_5_address0),
    .ce0(threshs_m_thresholds_5_ce0),
    .q0(threshs_m_thresholds_5_q0)
);

Thresholding_Batch_1_Thresholding_Batcg8j #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_4_address0),
    .ce0(threshs_m_thresholds_4_ce0),
    .q0(threshs_m_thresholds_4_q0)
);

Thresholding_Batch_1_Thresholding_Batchbi #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_3_address0),
    .ce0(threshs_m_thresholds_3_ce0),
    .q0(threshs_m_thresholds_3_q0)
);

Thresholding_Batch_1_Thresholding_Batcibs #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_2_address0),
    .ce0(threshs_m_thresholds_2_ce0),
    .q0(threshs_m_thresholds_2_q0)
);

Thresholding_Batch_1_Thresholding_BatcjbC #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_1_address0),
    .ce0(threshs_m_thresholds_1_ce0),
    .q0(threshs_m_thresholds_1_q0)
);

Thresholding_Batch_1_Thresholding_BatckbM #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_address0),
    .ce0(threshs_m_thresholds_ce0),
    .q0(threshs_m_thresholds_q0)
);

Thresholding_Batch_1_Thresholding_BatclbW #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_11_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_11_address0),
    .ce0(threshs_m_thresholds_11_ce0),
    .q0(threshs_m_thresholds_11_q0)
);

Thresholding_Batch_1_Thresholding_Batcmb6 #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_10_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_10_address0),
    .ce0(threshs_m_thresholds_10_ce0),
    .q0(threshs_m_thresholds_10_q0)
);

Thresholding_Batch_1_Thresholding_Batcncg #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_9_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_9_address0),
    .ce0(threshs_m_thresholds_9_ce0),
    .q0(threshs_m_thresholds_9_q0)
);

Thresholding_Batch_1_Thresholding_Batcocq #(
    .DataWidth( 19 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
threshs_m_thresholds_8_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(threshs_m_thresholds_8_address0),
    .ce0(threshs_m_thresholds_8_ce0),
    .q0(threshs_m_thresholds_8_q0)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_299_p2 == 1'd0))) begin
        i_0_reg_288 <= i_fu_305_p2;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_0_reg_288 <= 14'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_299_p2 == 1'd0))) begin
        nf_assign_reg_277 <= nf_1_fu_341_p3;
    end else if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        nf_assign_reg_277 <= 32'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        icmp_ln221_reg_720 <= icmp_ln221_fu_299_p2;
        icmp_ln221_reg_720_pp0_iter1_reg <= icmp_ln221_reg_720;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_reg_720 == 1'd0))) begin
        icmp_ln899_10_reg_872 <= icmp_ln899_10_fu_461_p2;
        icmp_ln899_11_reg_877 <= icmp_ln899_11_fu_470_p2;
        icmp_ln899_12_reg_882 <= icmp_ln899_12_fu_479_p2;
        icmp_ln899_13_reg_887 <= icmp_ln899_13_fu_488_p2;
        icmp_ln899_1_reg_827 <= icmp_ln899_1_fu_362_p2;
        icmp_ln899_2_reg_832 <= icmp_ln899_2_fu_371_p2;
        icmp_ln899_3_reg_837 <= icmp_ln899_3_fu_380_p2;
        icmp_ln899_4_reg_842 <= icmp_ln899_4_fu_389_p2;
        icmp_ln899_5_reg_847 <= icmp_ln899_5_fu_398_p2;
        icmp_ln899_6_reg_852 <= icmp_ln899_6_fu_407_p2;
        icmp_ln899_reg_822 <= icmp_ln899_fu_353_p2;
        xor_ln899_7_reg_857 <= xor_ln899_7_fu_421_p2;
        xor_ln899_8_reg_862 <= xor_ln899_8_fu_436_p2;
        xor_ln899_9_reg_867 <= xor_ln899_9_fu_451_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_299_p2 == 1'd0))) begin
        tmp_V_1_reg_729 <= in_V_V_TDATA;
    end
end

always @ (*) begin
    if ((icmp_ln221_fu_299_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state5) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state5)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln221_fu_299_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        in_V_V_TDATA_blk_n = in_V_V_TVALID;
    end else begin
        in_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_fu_299_p2 == 1'd0))) begin
        in_V_V_TREADY = 1'b1;
    end else begin
        in_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln221_reg_720_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        out_V_V_TDATA_blk_n = out_V_V_TREADY;
    end else begin
        out_V_V_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln221_reg_720_pp0_iter1_reg == 1'd0))) begin
        out_V_V_TVALID = 1'b1;
    end else begin
        out_V_V_TVALID = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_10_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_10_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_11_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_11_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_12_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_12_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_13_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_13_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_1_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_1_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_2_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_2_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_3_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_3_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_4_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_4_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_5_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_5_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_6_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_6_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_7_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_7_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_8_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_8_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_9_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_9_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        threshs_m_thresholds_ce0 = 1'b1;
    end else begin
        threshs_m_thresholds_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_299_p2 == 1'd1)) & ~((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_299_p2 == 1'd1)))) begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln700_10_fu_693_p2 = (zext_ln700_7_fu_689_p1 + zext_ln700_6_fu_679_p1);

assign add_ln700_11_fu_699_p2 = (add_ln700_10_fu_693_p2 + zext_ln700_5_fu_669_p1);

assign add_ln700_1_fu_615_p2 = (zext_ln700_1_fu_611_p1 + select_ln700_fu_498_p3);

assign add_ln700_2_fu_621_p2 = (zext_ln142_3_fu_529_p1 + zext_ln142_4_fu_538_p1);

assign add_ln700_3_fu_631_p2 = (zext_ln142_5_fu_547_p1 + zext_ln142_6_fu_556_p1);

assign add_ln700_4_fu_641_p2 = (zext_ln700_3_fu_637_p1 + zext_ln700_2_fu_627_p1);

assign add_ln700_5_fu_651_p2 = (zext_ln700_4_fu_647_p1 + add_ln700_1_fu_615_p2);

assign add_ln700_6_fu_657_p2 = (zext_ln142_8_fu_563_p1 + zext_ln142_9_fu_566_p1);

assign add_ln700_7_fu_663_p2 = (add_ln700_6_fu_657_p2 + zext_ln142_7_fu_560_p1);

assign add_ln700_8_fu_673_p2 = (zext_ln142_10_fu_574_p1 + zext_ln142_11_fu_583_p1);

assign add_ln700_9_fu_683_p2 = (zext_ln142_12_fu_592_p1 + zext_ln700_fu_601_p1);

assign add_ln700_fu_605_p2 = (zext_ln142_1_fu_511_p1 + zext_ln142_2_fu_520_p1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state5 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_299_p2 == 1'd0));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_block_state4_io)) | ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_299_p2 == 1'd0)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_block_state4_io)) | ((in_V_V_TVALID == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln221_fu_299_p2 == 1'd0)));
end

always @ (*) begin
    ap_block_state2_pp0_stage0_iter0 = ((in_V_V_TVALID == 1'b0) & (icmp_ln221_fu_299_p2 == 1'd0));
end

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state4_io = ((out_V_V_TREADY == 1'b0) & (icmp_ln221_reg_720_pp0_iter1_reg == 1'd0));
end

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign i_fu_305_p2 = (i_0_reg_288 + 14'd1);

assign icmp_ln221_fu_299_p2 = ((i_0_reg_288 == 14'd12800) ? 1'b1 : 1'b0);

assign icmp_ln235_fu_335_p2 = ((nf_fu_329_p2 == 32'd128) ? 1'b1 : 1'b0);

assign icmp_ln899_10_fu_461_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_10_fu_457_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_11_fu_470_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_11_fu_466_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_12_fu_479_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_12_fu_475_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_13_fu_488_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_13_fu_484_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_1_fu_362_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_1_fu_358_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_2_fu_371_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_2_fu_367_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_3_fu_380_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_3_fu_376_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_4_fu_389_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_4_fu_385_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_5_fu_398_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_5_fu_394_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_6_fu_407_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_6_fu_403_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_7_fu_416_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_7_fu_412_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_8_fu_431_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_8_fu_427_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_9_fu_446_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_9_fu_442_p1)) ? 1'b1 : 1'b0);

assign icmp_ln899_fu_353_p2 = (($signed(tmp_V_1_reg_729) < $signed(sext_ln142_fu_349_p1)) ? 1'b1 : 1'b0);

assign nf_1_fu_341_p3 = ((icmp_ln235_fu_335_p2[0:0] === 1'b1) ? 32'd0 : nf_fu_329_p2);

assign nf_fu_329_p2 = (nf_assign_reg_277 + 32'd1);

assign out_V_V_TDATA = tmp_V_fu_709_p2;

assign select_ln700_fu_498_p3 = ((xor_ln899_fu_493_p2[0:0] === 1'b1) ? 4'd10 : 4'd9);

assign sext_ln142_10_fu_457_p1 = $signed(threshs_m_thresholds_11_q0);

assign sext_ln142_11_fu_466_p1 = $signed(threshs_m_thresholds_10_q0);

assign sext_ln142_12_fu_475_p1 = $signed(threshs_m_thresholds_9_q0);

assign sext_ln142_13_fu_484_p1 = $signed(threshs_m_thresholds_8_q0);

assign sext_ln142_1_fu_358_p1 = $signed(threshs_m_thresholds_12_q0);

assign sext_ln142_2_fu_367_p1 = $signed(threshs_m_thresholds_7_q0);

assign sext_ln142_3_fu_376_p1 = $signed(threshs_m_thresholds_6_q0);

assign sext_ln142_4_fu_385_p1 = $signed(threshs_m_thresholds_5_q0);

assign sext_ln142_5_fu_394_p1 = $signed(threshs_m_thresholds_4_q0);

assign sext_ln142_6_fu_403_p1 = $signed(threshs_m_thresholds_3_q0);

assign sext_ln142_7_fu_412_p1 = $signed(threshs_m_thresholds_2_q0);

assign sext_ln142_8_fu_427_p1 = $signed(threshs_m_thresholds_1_q0);

assign sext_ln142_9_fu_442_p1 = $signed(threshs_m_thresholds_q0);

assign sext_ln142_fu_349_p1 = $signed(threshs_m_thresholds_13_q0);

assign threshs_m_thresholds_10_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_11_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_12_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_13_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_1_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_2_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_3_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_4_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_5_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_6_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_7_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_8_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_9_address0 = zext_ln142_fu_311_p1;

assign threshs_m_thresholds_address0 = zext_ln142_fu_311_p1;

assign tmp_V_fu_709_p2 = (zext_ln700_8_fu_705_p1 + add_ln700_5_fu_651_p2);

assign xor_ln899_10_fu_569_p2 = (icmp_ln899_10_reg_872 ^ 1'd1);

assign xor_ln899_11_fu_578_p2 = (icmp_ln899_11_reg_877 ^ 1'd1);

assign xor_ln899_12_fu_587_p2 = (icmp_ln899_12_reg_882 ^ 1'd1);

assign xor_ln899_13_fu_596_p2 = (icmp_ln899_13_reg_887 ^ 1'd1);

assign xor_ln899_1_fu_506_p2 = (icmp_ln899_1_reg_827 ^ 1'd1);

assign xor_ln899_2_fu_515_p2 = (icmp_ln899_2_reg_832 ^ 1'd1);

assign xor_ln899_3_fu_524_p2 = (icmp_ln899_3_reg_837 ^ 1'd1);

assign xor_ln899_4_fu_533_p2 = (icmp_ln899_4_reg_842 ^ 1'd1);

assign xor_ln899_5_fu_542_p2 = (icmp_ln899_5_reg_847 ^ 1'd1);

assign xor_ln899_6_fu_551_p2 = (icmp_ln899_6_reg_852 ^ 1'd1);

assign xor_ln899_7_fu_421_p2 = (icmp_ln899_7_fu_416_p2 ^ 1'd1);

assign xor_ln899_8_fu_436_p2 = (icmp_ln899_8_fu_431_p2 ^ 1'd1);

assign xor_ln899_9_fu_451_p2 = (icmp_ln899_9_fu_446_p2 ^ 1'd1);

assign xor_ln899_fu_493_p2 = (icmp_ln899_reg_822 ^ 1'd1);

assign zext_ln142_10_fu_574_p1 = xor_ln899_10_fu_569_p2;

assign zext_ln142_11_fu_583_p1 = xor_ln899_11_fu_578_p2;

assign zext_ln142_12_fu_592_p1 = xor_ln899_12_fu_587_p2;

assign zext_ln142_1_fu_511_p1 = xor_ln899_1_fu_506_p2;

assign zext_ln142_2_fu_520_p1 = xor_ln899_2_fu_515_p2;

assign zext_ln142_3_fu_529_p1 = xor_ln899_3_fu_524_p2;

assign zext_ln142_4_fu_538_p1 = xor_ln899_4_fu_533_p2;

assign zext_ln142_5_fu_547_p1 = xor_ln899_5_fu_542_p2;

assign zext_ln142_6_fu_556_p1 = xor_ln899_6_fu_551_p2;

assign zext_ln142_7_fu_560_p1 = xor_ln899_7_reg_857;

assign zext_ln142_8_fu_563_p1 = xor_ln899_8_reg_862;

assign zext_ln142_9_fu_566_p1 = xor_ln899_9_reg_867;

assign zext_ln142_fu_311_p1 = nf_assign_reg_277;

assign zext_ln700_1_fu_611_p1 = add_ln700_fu_605_p2;

assign zext_ln700_2_fu_627_p1 = add_ln700_2_fu_621_p2;

assign zext_ln700_3_fu_637_p1 = add_ln700_3_fu_631_p2;

assign zext_ln700_4_fu_647_p1 = add_ln700_4_fu_641_p2;

assign zext_ln700_5_fu_669_p1 = add_ln700_7_fu_663_p2;

assign zext_ln700_6_fu_679_p1 = add_ln700_8_fu_673_p2;

assign zext_ln700_7_fu_689_p1 = add_ln700_9_fu_683_p2;

assign zext_ln700_8_fu_705_p1 = add_ln700_11_fu_699_p2;

assign zext_ln700_fu_601_p1 = xor_ln899_13_fu_596_p2;

endmodule //Thresholding_Batch_1_Thresholding_Batch
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActEe0.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActEe0_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActEe0_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActEe0(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActEe0_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActEe0_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActBew.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActBew_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActBew_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActBew(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActBew_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActBew_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbFp.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcbFp_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbFp_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcbFp(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcbFp_rom Thresholding_Batch_0_Thresholding_BatcbFp_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActAem.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActAem_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 18;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActAem_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActAem(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd18;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActAem_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActAem_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actzec.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Actzec_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Actzec_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Actzec(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Actzec_rom StreamingFCLayer_Batch_2_Matrix_Vector_Actzec_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/e911/Q_srl.v

// original source:
// https://github.com/nachiket/tdfc/blob/master/verilog/queues/Q_srl_oreg3_prefull_SIMPLE.v


// Copyright (c) 1999 The Regents of the University of California
// Copyright (c) 2010 The Regents of the University of Pennsylvania
// Copyright (c) 2011 Department of Electrical and Electronic Engineering, Imperial College London
// Copyright (c) 2020 Xilinx
//
// Permission to use, copy, modify, and distribute this software and
// its documentation for any purpose, without fee, and without a
// written agreement is hereby granted, provided that the above copyright
// notice and this paragraph and the following two paragraphs appear in
// all copies.
//
// IN NO EVENT SHALL THE UNIVERSITY OF CALIFORNIA BE LIABLE TO ANY PARTY FOR
// DIRECT, INDIRECT, SPECIAL, INCIDENTAL, OR CONSEQUENTIAL DAMAGES, INCLUDING
// LOST PROFITS, ARISING OUT OF THE USE OF THIS SOFTWARE AND ITS DOCUMENTATION,
// EVEN IF THE UNIVERSITY OF CALIFORNIA HAS BEEN ADVISED OF THE POSSIBILITY OF
// SUCH DAMAGE.
//
// THE UNIVERSITY OF CALIFORNIA SPECIFICALLY DISCLAIMS ANY WARRANTIES,
// INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
// AND FITNESS FOR A PARTICULAR PURPOSE. THE SOFTWARE PROVIDED HEREUNDER IS ON
// AN "AS IS" BASIS, AND THE UNIVERSITY OF CALIFORNIA HAS NO OBLIGATIONS TO
// PROVIDE MAINTENANCE, SUPPORT, UPDATES, ENHANCEMENTS, OR MODIFICATIONS.
//

// Q_srl_oreg3_prefull_SIMPLE.v
//
//  - In-page queue with parameterizable depth, bit width
//  - Stream I/O is triple (data, valid, back-pressure),
//      with EOS concatenated into the data
//  - Flow control for input & output is combinationally decoupled
//  - 2 <= depth <= 256
//      * (depth >= 2)  is required to decouple I/O flow control,
//          where empty => no produce,  full => no consume,
//          and depth 1 would ping-pong between the two at half rate
//      * (depth <= 256) can be modified
//           by changing ''synthesis loop_limit X'' below
//          and changing ''addrwidth'' or its log computation
//  - 1 <= width
//  - Queue storage is in SRL16E, up to depth 16 per LUT per bit-slice,
//      plus output register (for fast output)
//  - Queue addressing is done by ''addr'' up-down counter
//  - Queue fullness is checked by comparator (addr==depth)
//  - Queue fullness                           is pre-computed for next cycle
//  - Queue input back-pressure                is pre-computed for next cycle
//  - Queue output valid (state!=state__empty) is pre-computed for next cycle
//      (necessary since SRL data output reg requires non-boolean state)
//  - FSM has 3 states (empty, one, more)
//  - When empty, continue to emit most recently emitted value (for debugging)
//
//  - Queue slots used      = / (state==state_empty) ? 0
//                            | (state==state_one)   ? 1
//                            \ (state==state_more)  ? addr+2
//  - Queue slots used     <=  depth
//  - Queue slots remaining =  depth - used
//                          = / (state==state_empty) ? depth
//                            | (state==state_one)   ? depth-1
//                            \ (state==state_more)  ? depth-2-addr
//
//  - Synplify 7.1 / 8.0
//  - Eylon Caspi,  9/11/03, 8/18/04, 3/29/05


`ifdef  Q_srl
`else
`define Q_srl


module Q_srl (clock, reset, i_d, i_v, i_r, o_d, o_v, o_r, count);

   parameter depth = 16;   // - greatest #items in queue  (2 <= depth <= 256)
   parameter width = 16;   // - width of data (i_d, o_d)

   parameter addrwidth = $clog2(depth);

   input     clock;
   input     reset;

   input  [width-1:0] i_d;	// - input  stream data (concat data + eos)
   input              i_v;	// - input  stream valid
   output             i_r;	// - input  stream ready
   wire               i_b;  // - input  stream back-pressure

   output [width-1:0] o_d;	// - output stream data (concat data + eos)
   output             o_v;	// - output stream valid
   input              o_r;	// - output stream ready
   wire               o_b;	// - output stream back-pressure

   output [addrwidth:0] count;  // - output number of elems in queue

   reg    [addrwidth-1:0] addr, addr_, a_;		// - SRL16 address
							//     for data output
   reg 			  shift_en_;			// - SRL16 shift enable
   reg    [width-1:0] 	  srl [depth-2:0];		// - SRL16 memory
   reg 			  shift_en_o_;			// - SRLO  shift enable
   reg    [width-1:0] 	  srlo_, srlo			// - SRLO  output reg
			  /* synthesis syn_allow_retiming=0 */ ;

   parameter state_empty = 2'd0;    // - state empty : o_v=0 o_d=UNDEFINED
   parameter state_one   = 2'd1;    // - state one   : o_v=1 o_d=srlo
   parameter state_more  = 2'd2;    // - state more  : o_v=1 o_d=srlo
				    //     #items in srl = addr+2

   reg [1:0] state, state_;	    // - state register

   wire      addr_full_;	    // - true iff addr==depth-2 on NEXT cycle
   reg       addr_full; 	    // - true iff addr==depth-2
   wire      addr_zero_;	    // - true iff addr==0
   wire      o_v_reg_;		    // - true iff state_empty   on NEXT cycle
   reg       o_v_reg  		    // - true iff state_empty
	     /* synthesis syn_allow_retiming=0 */ ;
   wire      i_b_reg_;		    // - true iff !full         on NEXT cycle
   reg       i_b_reg  		    // - true iff !full
	     /* synthesis syn_allow_retiming=0 */ ;

   assign addr_full_ = (state_==state_more) && (addr_==depth-2);
						// - queue full
   assign addr_zero_ = (addr==0);		// - queue contains 2 (or 1,0)
   assign o_v_reg_   = (state_!=state_empty);	// - output valid if non-empty
   assign i_b_reg_   = addr_full_;		// - input bp if full
   assign o_d = srlo;				// - output data from queue
   assign o_v = o_v_reg;			// - output valid if non-empty
   assign i_b = i_b_reg;			// - input bp if full

   assign i_r = !i_b;
   assign o_b = !o_r;

   assign count = (state==state_more ? addr+2 : (state==state_one ? 1 : 0));

   // - ''always'' block with both FFs and SRL16 does not work,
   //      since FFs need reset but SRL16 does not

   always @(posedge clock) begin	// - seq always: FFs
      if (reset) begin
	 state     <= state_empty;
	 addr      <= 0;
         addr_full <= 0;
	 o_v_reg   <= 0;
	 i_b_reg   <= 1;
      end
      else begin
	 state     <= state_;
	 addr      <= addr_;
         addr_full <= addr_full_;
	 o_v_reg   <= o_v_reg_;
	 i_b_reg   <= i_b_reg_;
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin	// - seq always: srlo
      // - infer enabled output reg at end of shift chain
      // - input first element from i_d, all subsequent elements from SRL16
      if (reset) begin
	 srlo <= 0;
      end
      else begin
	 if (shift_en_o_) begin
	    srlo <= srlo_;
	 end
      end
   end // always @ (posedge clock)

   always @(posedge clock) begin			// - seq always: srl
      // - infer enabled SRL16E from shifting srl array
      // - no reset capability;  srl[] contents undefined on reset
      if (shift_en_) begin
	 // synthesis loop_limit 256
	 for (a_=depth-2; a_>0; a_=a_-1) begin
	    srl[a_] = srl[a_-1];
	 end
	 srl[0] <= i_d;
      end
   end // always @ (posedge clock or negedge reset)

   always @* begin					// - combi always
        srlo_       <=  'bx;
        shift_en_o_ <= 1'bx;
        shift_en_   <= 1'bx;
        addr_       <=  'bx;
        state_      <= 2'bx;
      case (state)

	state_empty: begin		    // - (empty, will not produce)
	      if (i_v) begin		    // - empty & i_v => consume
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else	begin		    // - empty & !i_v => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end

	state_one: begin		    // - (contains one)
	      if (i_v && o_b) begin	    // - one & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - one & i_v & !o_b => cons+prod
		 srlo_       <= i_d;
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && o_b) begin   // - one & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_one;
	      end
	      else if (!i_v && !o_b) begin  // - one & !i_v & !o_b => produce
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1'bx;
		 addr_       <= 0;
		 state_      <= state_empty;
	      end
	end // case: state_one

	state_more: begin		    // - (contains more than one)
	   if (addr_full || (depth==2)) begin
					    // - (full, will not consume)
					    // - (full here if depth==2)
	      if (o_b) begin		    // - full & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else begin		    // - full & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
//		 addr_       <= addr-1;
//		 state_      <= state_more;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end
	   else begin			    // - (mid: neither empty nor full)
	      if (i_v && o_b) begin	    // - mid & i_v & o_b => consume
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 1;
		 addr_       <= addr+1;
		 state_      <= state_more;
	      end
	      else if (i_v && !o_b) begin   // - mid & i_v & !o_b => cons+prod
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 1;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && o_b) begin   // - mid & !i_v & o_b => idle
		 srlo_       <= 'bx;
		 shift_en_o_ <= 0;
		 shift_en_   <= 0;
		 addr_       <= addr;
		 state_      <= state_more;
	      end
	      else if (!i_v && !o_b) begin  // - mid & !i_v & !o_b => produce
		 srlo_       <= srl[addr];
		 shift_en_o_ <= 1;
		 shift_en_   <= 0;
		 addr_       <= addr_zero_ ? 0         : addr-1;
		 state_      <= addr_zero_ ? state_one : state_more;
	      end
	   end // else: !if(addr_full)
	end // case: state_more

	default: begin
		 srlo_       <=  'bx;
		 shift_en_o_ <= 1'bx;
		 shift_en_   <= 1'bx;
		 addr_       <=  'bx;
		 state_      <= 2'bx;
	end // case: default

      endcase // case(state)
   end // always @ *

endmodule // Q_srl


`endif  // `ifdef  Q_srl
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcbkb.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_Batcbkb_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_Batcbkb_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_Batcbkb(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_Batcbkb_rom Thresholding_Batch_1_Thresholding_Batcbkb_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccGz.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatccGz_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 8;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatccGz_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatccGz(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd8;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatccGz_rom Thresholding_Batch_0_Thresholding_BatccGz_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcNgs.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcNgs_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcNgs_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcNgs(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcNgs_rom Thresholding_Batch_0_Thresholding_BatcNgs_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/6e26/StreamingFIFO_18.v


module StreamingFIFO_18(
ap_clk,
ap_rst_n,
count,
in0_V_V_TDATA,
in0_V_V_TVALID,
in0_V_V_TREADY,
out_V_V_TDATA,
out_V_V_TVALID,
out_V_V_TREADY
);

input   ap_clk;
input   ap_rst_n;
output [13:0] count;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [15:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

Q_srl #(
.depth(16384),
.width(16)
)
StreamingFIFO_18_StreamingFIFO_18
(
 .clock(ap_clk),
 .reset(!ap_rst_n),
 .count(count),
 .i_d(in0_V_V_TDATA),
 .i_v(in0_V_V_TVALID),
 .i_r(in0_V_V_TREADY),
 .o_d(out_V_V_TDATA),
 .o_v(out_V_V_TVALID),
 .o_r(out_V_V_TREADY)
);

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcjbC.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcjbC_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 4;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcjbC_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcjbC(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd4;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcjbC_rom Thresholding_Batch_0_Thresholding_BatcjbC_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/a3f1/hdl/verilog/ConvolutionInputGenerator_1_ConvolutionInputGfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module ConvolutionInputGenerator_1_ConvolutionInputGfYi #(
parameter
    ID                = 0,
    NUM_STAGE         = 1,
    din0_WIDTH       = 32,
    din1_WIDTH       = 32,
    din2_WIDTH       = 32,
    din3_WIDTH       = 32,
    din4_WIDTH         = 32,
    dout_WIDTH            = 32
)(
    input  [15 : 0]     din0,
    input  [15 : 0]     din1,
    input  [15 : 0]     din2,
    input  [15 : 0]     din3,
    input  [1 : 0]    din4,
    output [15 : 0]   dout);

// puts internal signals
wire [1 : 0]     sel;
// level 1 signals
wire [15 : 0]         mux_1_0;
wire [15 : 0]         mux_1_1;
// level 2 signals
wire [15 : 0]         mux_2_0;

assign sel = din4;

// Generate level 1 logic
assign mux_1_0 = (sel[0] == 0)? din0 : din1;
assign mux_1_1 = (sel[0] == 0)? din2 : din3;

// Generate level 2 logic
assign mux_2_0 = (sel[1] == 0)? mux_1_0 : mux_1_1;

// output logic
assign dout = mux_2_0;

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbDo.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcbDo_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcbDo_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcbDo(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcbDo_rom Thresholding_Batch_0_Thresholding_BatcbDo_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActJfO.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActJfO_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActJfO_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActJfO(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActJfO_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActJfO_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcThq.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcThq_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 6;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcThq_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcThq(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd6;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcThq_rom Thresholding_Batch_0_Thresholding_BatcThq_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0da3/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActDeQ.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActDeQ_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_3_u6fssgdv/project_StreamingFCLayer_Batch_3/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_3_Matrix_Vector_ActDeQ_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_3_Matrix_Vector_ActDeQ(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_3_Matrix_Vector_ActDeQ_rom StreamingFCLayer_Batch_3_Matrix_Vector_ActDeQ_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/3a3d/hdl/verilog/StreamingDataWidthConverter_Batch_2_StreamingDataWidthConverter_Batch_2.v

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2020.1.1
// Copyright (C) 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="StreamingDataWidthConverter_Batch_2_StreamingDataWidthConverter_Batch_2,hls_ip_2020_1_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=1,HLS_INPUT_PART=xc7z020-clg400-1,HLS_INPUT_CLOCK=10.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=5.025000,HLS_SYN_LAT=69,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=115,HLS_SYN_LUT=223,HLS_VERSION=2020_1_1}" *)

module StreamingDataWidthConverter_Batch_2_StreamingDataWidthConverter_Batch_2 (
        ap_clk,
        ap_rst_n,
        in0_V_V_TDATA,
        in0_V_V_TVALID,
        in0_V_V_TREADY,
        out_V_V_TDATA,
        out_V_V_TVALID,
        out_V_V_TREADY
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst_n;
input  [15:0] in0_V_V_TDATA;
input   in0_V_V_TVALID;
output   in0_V_V_TREADY;
output  [31:0] out_V_V_TDATA;
output   out_V_V_TVALID;
input   out_V_V_TREADY;

reg in0_V_V_TREADY;

 reg    ap_rst_n_inv;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_start;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_done;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_idle;
wire    grp_StreamingDataWidthCo_1_fu_26_ap_ready;
wire    grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
wire   [31:0] grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID;
wire    grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY;
reg    grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;
(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
reg   [3:0] ap_NS_fsm;
wire    ap_CS_fsm_state4;
wire    regslice_both_out_V_V_U_apdone_blk;
wire    regslice_both_in0_V_V_U_apdone_blk;
wire   [15:0] in0_V_V_TDATA_int;
wire    in0_V_V_TVALID_int;
reg    in0_V_V_TREADY_int;
wire    regslice_both_in0_V_V_U_ack_in;
wire    out_V_V_TREADY_int;
wire    regslice_both_out_V_V_U_vld_out;

// power-on initialization
initial begin
#0 grp_StreamingDataWidthCo_1_fu_26_ap_start_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
end

StreamingDataWidthConverter_Batch_2_StreamingDataWidthCo_1 grp_StreamingDataWidthCo_1_fu_26(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_StreamingDataWidthCo_1_fu_26_ap_start),
    .ap_done(grp_StreamingDataWidthCo_1_fu_26_ap_done),
    .ap_idle(grp_StreamingDataWidthCo_1_fu_26_ap_idle),
    .ap_ready(grp_StreamingDataWidthCo_1_fu_26_ap_ready),
    .in_V_V_TDATA(in0_V_V_TDATA_int),
    .in_V_V_TVALID(in0_V_V_TVALID_int),
    .in_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY),
    .out_V_V_TDATA(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .out_V_V_TVALID(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .out_V_V_TREADY(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY)
);

regslice_both #(
    .DataWidth( 16 ))
regslice_both_in0_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(in0_V_V_TDATA),
    .vld_in(in0_V_V_TVALID),
    .ack_in(regslice_both_in0_V_V_U_ack_in),
    .data_out(in0_V_V_TDATA_int),
    .vld_out(in0_V_V_TVALID_int),
    .ack_out(in0_V_V_TREADY_int),
    .apdone_blk(regslice_both_in0_V_V_U_apdone_blk)
);

regslice_both #(
    .DataWidth( 32 ))
regslice_both_out_V_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TDATA),
    .vld_in(grp_StreamingDataWidthCo_1_fu_26_out_V_V_TVALID),
    .ack_in(out_V_V_TREADY_int),
    .data_out(out_V_V_TDATA),
    .vld_out(regslice_both_out_V_V_U_vld_out),
    .ack_out(out_V_V_TREADY),
    .apdone_blk(regslice_both_out_V_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b1;
        end else if ((grp_StreamingDataWidthCo_1_fu_26_ap_ready == 1'b1)) begin
            grp_StreamingDataWidthCo_1_fu_26_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_in0_V_V_U_ack_in == 1'b1) & (in0_V_V_TVALID == 1'b1))) begin
        in0_V_V_TREADY = 1'b1;
    end else begin
        in0_V_V_TREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        in0_V_V_TREADY_int = grp_StreamingDataWidthCo_1_fu_26_in_V_V_TREADY;
    end else begin
        in0_V_V_TREADY_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            if (((grp_StreamingDataWidthCo_1_fu_26_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((regslice_both_out_V_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign grp_StreamingDataWidthCo_1_fu_26_ap_start = grp_StreamingDataWidthCo_1_fu_26_ap_start_reg;

assign grp_StreamingDataWidthCo_1_fu_26_out_V_V_TREADY = (out_V_V_TREADY_int & ap_CS_fsm_state3);

assign out_V_V_TVALID = regslice_both_out_V_V_U_vld_out;

endmodule //StreamingDataWidthConverter_Batch_2_StreamingDataWidthConverter_Batch_2
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcwdI.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_BatcwdI_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 5;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_BatcwdI_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_BatcwdI(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd5;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_BatcwdI_rom Thresholding_Batch_0_Thresholding_BatcwdI_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/209a/hdl/axilite_if.v

/*
 Copyright (c) 2020, Xilinx
 All rights reserved.

 Redistribution and use in source and binary forms, with or without
 modification, are permitted provided that the following conditions are met:

 * Redistributions of source code must retain the above copyright notice, this
   list of conditions and the following disclaimer.

 * Redistributions in binary form must reproduce the above copyright notice,
   this list of conditions and the following disclaimer in the documentation
   and/or other materials provided with the distribution.

 * Neither the name of FINN nor the names of its
   contributors may be used to endorse or promote products derived from
   this software without specific prior written permission.

 THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
 FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
 SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
 CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
 OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

module axi4lite_if
#(
    parameter ADDR_WIDTH = 32,
    parameter DATA_WIDTH = 32,//AXI4 spec requires this to be strictly 32 or 64
    parameter IP_DATA_WIDTH = 64//can be any power-of-2 multiple of DATA_WIDTH
)
(
//system signals
input aclk,
input aresetn,//active low, asynchronous assertion and synchronous deassertion

//Write channels
//write address
output reg                  awready,
input                       awvalid,
input [ADDR_WIDTH-1:0]      awaddr,
input [2:0]                 awprot,
//write data
output reg                  wready,
input                       wvalid,
input [DATA_WIDTH-1:0]      wdata,
input [(DATA_WIDTH/8)-1:0]  wstrb,
//burst response
input                       bready,
output reg                  bvalid,
output reg [1:0]            bresp,//NOTE: 00 = OKAY, 10 = SLVERR (write error)

//Read channels
//read address
output reg                  arready,
input                       arvalid,
input [ADDR_WIDTH-1:0]      araddr,
input [2:0]                 arprot,
//read data
input                       rready,
output reg                  rvalid,
output reg [1:0]            rresp,//NOTE: 00 = OKAY, 10 = SLVERR (read error)
output reg [DATA_WIDTH-1:0] rdata,

//IP-side interface
output reg                  ip_en,
output reg                  ip_wen,
output reg [ADDR_WIDTH-1:0] ip_addr,
output [IP_DATA_WIDTH-1:0]  ip_wdata,
input                       ip_rack,
input [IP_DATA_WIDTH-1:0]      ip_rdata
);

localparam RESP_OKAY = 2'b00;
localparam RESP_SLVERR = 2'b10;
//get ceil(log2(ceil(IP_DATA_WIDTH/DATA_WIDTH)))
localparam NFOLDS_LOG = $clog2((IP_DATA_WIDTH + DATA_WIDTH - 1) / DATA_WIDTH);

reg                      internal_ren;
reg                      internal_wen;
reg                      internal_wack;
reg [ADDR_WIDTH-1:0]     internal_raddr;
reg [ADDR_WIDTH-1:0]     internal_waddr;
reg [DATA_WIDTH-1:0]     internal_wdata;
wire [DATA_WIDTH-1:0]    internal_rdata;
reg                      internal_error = 0;

//check DATA_WIDTH
initial begin
    if(DATA_WIDTH != 32 & DATA_WIDTH != 64) begin
        $display("AXI4Lite DATA_WIDTH must be 32 or 64");
        $finish;
    end
end

//transaction state machine
localparam  STATE_IDLE  = 0,
            STATE_READ  = 1,
            STATE_WRITE = 2;

reg [1:0] state;

always @(posedge aclk or negedge aresetn)
    if(~aresetn)
        state <= STATE_IDLE;
    else case(state)
        STATE_IDLE:
            if(awvalid & wvalid)
                state <= STATE_WRITE;
            else if(arvalid)
                state <= STATE_READ;
        STATE_READ:
            if(rvalid & rready)
                state <= STATE_IDLE;
        STATE_WRITE:
            if(bvalid & bready)
                state <= STATE_IDLE;
        default: state <= STATE_IDLE;
    endcase

//write-related internal signals
always @(*) begin
    internal_waddr = awaddr >> $clog2(DATA_WIDTH/8);
    internal_wdata = wdata;
    internal_wen = (state == STATE_IDLE) & awvalid & wvalid;
end

always @(posedge aclk) begin
    awready <= internal_wen;
    wready <= internal_wen;
end

//read-related internal signals
always @(*) begin
    internal_raddr = araddr >> $clog2(DATA_WIDTH/8);
    internal_ren = (state == STATE_IDLE) & ~internal_wen & arvalid;
end

always @(posedge aclk)
    arready <= internal_ren;

wire write_to_last_fold;

always @(posedge aclk) begin
    ip_wen <= write_to_last_fold;
    ip_en <= internal_ren | write_to_last_fold;
    if(internal_ren | write_to_last_fold)
        ip_addr <= internal_ren ? (internal_raddr >> NFOLDS_LOG) : (internal_waddr >> NFOLDS_LOG);
    internal_wack <= internal_wen;
end

genvar i;
reg [(1<<NFOLDS_LOG)*DATA_WIDTH-1:0] ip_wdata_wide;
generate
if(NFOLDS_LOG == 0) begin: no_fold
    assign write_to_last_fold = internal_wen;
    assign internal_rdata = ip_rdata;
    always @(posedge aclk)
        ip_wdata_wide <= internal_wdata;
end else begin: fold
    reg [NFOLDS_LOG-1:0] internal_rfold;
    assign write_to_last_fold = internal_wen & (internal_waddr[NFOLDS_LOG-1:0] == {(NFOLDS_LOG){1'b1}});
    assign internal_rdata = ip_rdata >> (internal_rfold*DATA_WIDTH);
    always @(posedge aclk)
        if(internal_ren)
            internal_rfold <= internal_raddr[NFOLDS_LOG-1:0];
    for(i=0; i<(1<<NFOLDS_LOG); i = i+1) begin: gen_wdata
        always @(posedge aclk)
            if(internal_waddr[NFOLDS_LOG-1:0] == i)
                ip_wdata_wide[(i+1)*DATA_WIDTH-1:i*DATA_WIDTH] <= internal_wdata;
    end
end
endgenerate
assign ip_wdata = ip_wdata_wide[IP_DATA_WIDTH-1:0];

//write response on AXI4L bus
always @(posedge aclk or negedge aresetn)
    if(~aresetn) begin
        bvalid <= 0;//AXI4 spec requires BVALID pulled LOW during reset
        bresp <= RESP_OKAY;
    end else if(internal_wack) begin
        bvalid <= 1;
        bresp <= internal_error ? RESP_SLVERR : RESP_OKAY;
    end else if(bready) begin
        bvalid <= 0;
        bresp <= RESP_OKAY;
    end

//read response on AXI4L bus
always @(posedge aclk or negedge aresetn)
    if(~aresetn) begin
        rvalid <= 0;//AXI4 spec requires RVALID pulled LOW during reset
        rdata <= 0;
        rresp <= RESP_OKAY;
    end else if(ip_rack) begin
        rvalid <= 1;
        rdata <= internal_rdata;
        rresp <= internal_error ? RESP_SLVERR : RESP_OKAY;
    end else if(rready) begin
        rvalid <= 0;
        rdata <= 0;
        rresp <= RESP_OKAY;
    end

endmodule
//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/8864/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Acttde.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module StreamingFCLayer_Batch_2_Matrix_Vector_Acttde_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_2_4yckv8t4/project_StreamingFCLayer_Batch_2/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_2_Matrix_Vector_Acttde_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_2_Matrix_Vector_Acttde(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_2_Matrix_Vector_Acttde_rom StreamingFCLayer_Batch_2_Matrix_Vector_Acttde_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActZio.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActZio_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActZio_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActZio(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActZio_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActZio_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActfYi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActfYi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActfYi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActfYi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActfYi_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActfYi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/0fa4/hdl/verilog/Thresholding_Batch_1_Thresholding_Batchbi.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_1_Thresholding_Batchbi_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 19;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_1_wv2afg1v/project_Thresholding_Batch_1/sol1/impl/ip/hdl/verilog/Thresholding_Batch_1_Thresholding_Batchbi_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_1_Thresholding_Batchbi(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd19;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_1_Thresholding_Batchbi_rom Thresholding_Batch_1_Thresholding_Batchbi_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActFfa.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActFfa_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActFfa_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActFfa(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActFfa_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActFfa_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4ac7/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbrm.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module Thresholding_Batch_0_Thresholding_Batcbrm_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 7;
parameter AWIDTH = 2;
parameter MEM_SIZE = 3;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

(* ram_style = "distributed" *)reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_Thresholding_Batch_0_3w_u_csh/project_Thresholding_Batch_0/sol1/impl/ip/hdl/verilog/Thresholding_Batch_0_Thresholding_Batcbrm_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module Thresholding_Batch_0_Thresholding_Batcbrm(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd7;
parameter AddressRange = 32'd3;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



Thresholding_Batch_0_Thresholding_Batcbrm_rom Thresholding_Batch_0_Thresholding_Batcbrm_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/4b6a/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActlbW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActlbW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_4_2kaxius9/project_StreamingFCLayer_Batch_4/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_4_Matrix_Vector_ActlbW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_4_Matrix_Vector_ActlbW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_4_Matrix_Vector_ActlbW_rom StreamingFCLayer_Batch_4_Matrix_Vector_ActlbW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

//Added from /home/grgov/Diplomski_rad/finn_modified_docker_output_dir/vivado_stitch_proj_db1z4qol/finn_vivado_stitch_proj.srcs/sources_1/bd/finn_design/ipshared/156f/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActQgW.v

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2020.1.1 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActQgW_rom (
addr0, ce0, q0, clk);

parameter DWIDTH = 17;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output reg[DWIDTH-1:0] q0;
input clk;

reg [DWIDTH-1:0] ram[0:MEM_SIZE-1];

initial begin
    $readmemh("/home/grgov/Diplomski_rad/finn_modified_docker_output_dir/code_gen_ipgen_StreamingFCLayer_Batch_1_gj26dggu/project_StreamingFCLayer_Batch_1/sol1/impl/ip/hdl/verilog/StreamingFCLayer_Batch_1_Matrix_Vector_ActQgW_rom.dat", ram);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram[addr0];
    end
end



endmodule

`timescale 1 ns / 1 ps
module StreamingFCLayer_Batch_1_Matrix_Vector_ActQgW(
    reset,
    clk,
    address0,
    ce0,
    q0);

parameter DataWidth = 32'd17;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;



StreamingFCLayer_Batch_1_Matrix_Vector_ActQgW_rom StreamingFCLayer_Batch_1_Matrix_Vector_ActQgW_rom_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ));

endmodule

